//////////////////////////////////////////////////////////////////////
// JVS Controller Module for Analogizer - ALPHA VERSION
// Partial JVS Master implementation optimized for gaming performance
// 
// ⚠️  ALPHA STATUS - PARTIAL COMMAND IMPLEMENTATION ⚠️
//
// This module implements a JVS (JAMMA Video Standard) Master controller
// that allows connecting JVS arcade cabinets to the Analogue Pocket 
// through the Analogizer.
//
// IMPLEMENTATION STATUS (ALPHA ~30-40% complete):
// Based on JVS Specification v3.0 (25 pages, 49 commands total)
//
// ✅ FULLY IMPLEMENTED (8/49 commands):
//    - Reset (F0) - Double reset sequence with timing delays
//    - Set Address (F1) - Single device addressing
//    - IO Identity (10) - Device name string reading (up to 100 chars)
//    - Command Revision (11) - Format revision detection (BCD)
//    - JVS Revision (12) - Protocol version detection (BCD) 
//    - Communications Version (13) - Communication system version
//    - Feature Check (14) - Complete capability parsing with all function codes
//    - Switch Inputs (20) - Digital buttons (2 players, 13 buttons each)
//    - Analog Inputs (22) - Multi-channel 16-bit analog data
//    - Generic Output 1 (32) - Digital GPIO control (3-byte format)
//    - JVS escape sequences (D0 DF → E0, D0 CF → D0)
//    - RS485 timing control with setup/hold delays
//
// 🟡 PARTIALLY IMPLEMENTED (4/49 commands):
//    - Coin Inputs (21) - Command sent, status parsed but coin data ignored
//    - Screen Position Inputs (25) - Basic X/Y coordinates (16-bit each)
//    - Keycode Inputs (24) - Command sent, response skipped
//    - Misc Switch Inputs (26) - Command sent, response skipped
//
// ❌ NOT IMPLEMENTED (37/49 commands):
//    - Main ID (15) - Send main board identification to device
//    - Rotary Inputs (23) - Rotary encoder data (parsed but ignored)
//    - Remaining Payout (2E) - Medal hopper status and count
//    - Data Retransmit (2F) - Checksum error recovery
//    - Coin management: COINDEC (30), COININC (35), PAYINC (31), PAYDEC (36)
//    - Advanced outputs: OUTPUT2 (37), OUTPUT3 (38), ANLOUT (33), CHAROUT (34)
//    - Communication changes: COMMCHG (F2)
//    - Manufacturer-specific commands (Taito TypeX, Namco, CyberLead LED)
//    - Multi-device addressing (supports single device only)
//    - Dynamic baud rate changes
//    - Error recovery mechanisms
//
// PLANNED RESTRUCTURING:
// This monolithic module will be split into:
//   - jvs_com: Communication layer (UART, framing, escape sequences)
//   - jvs_controller: Protocol layer (commands, parsing, state machines)
//   - SNAC interface abstraction: Review interaction with SNAC module for
//     better abstraction and future portability to MiSTer platform
//
// ARCHITECTURE (Current):
// - RS485 State Machine: Manages transceiver direction and timing
// - Main State Machine: Handles JVS protocol sequence and commands  
// - RX State Machine: Processes incoming JVS responses with full parsing
// - Two-buffer system: Raw buffer + processed buffer for unescaped data
// - Node information management for device capabilities
//
// PROTOCOL COMPLIANCE:
// - Physical Layer: RS-485 at 115200 baud (8N1) ✅
// - Link Layer: SYNC(0xE0) + NODE + LENGTH + DATA + CHECKSUM ✅  
// - Escape sequences: D0 DF → E0, D0 CF → D0 ✅
// - Address assignment: Master=0x00, Slaves=0x01-0x1F ✅
// - Initialization: Double reset + sequential addressing ✅
// - Multi-device chaining: Infrastructure present but single device only
//
// HARDWARE REQUIREMENTS:
// - External MAX485 or equivalent RS485 transceiver
// - Proper 120Ω termination for reliable communication  
// - JVS-compatible arcade cabinet
// - SENSE line connection for proper device chaining (unused in single mode)
//
// I/O BOARD COMPATIBILITY:
// ✅ WORKING:
//    - NAJV2 (Tekken 7) - Full compatibility
//    - NAJV (Time Crisis 4) - Full compatibility  
//    - TAITO CORP Ver2.0 (Viewlix) - Full compatibility
// ❌ NOT WORKING:
//    - "No Brand;NAOMI Converter98701;ver2.0" - Frames ignored
//
// Author: Totaly FuRy - Sebastien DUPONCHEEL (sduponch on GitHub)
// Project: Analogizer JVS Controller
// Status: Alpha - Partial Implementation
// Date: 2025
//////////////////////////////////////////////////////////////////////
//Use: set_global_assignment -name VERILOG_MACRO "USE_DUMMY_JVS_DATA=1" 
//in project .qsf to use dummy data for simulation without JVS device

`default_nettype none
`timescale 1ns / 1ps

import jvs_node_info_pkg::*;

module jvs_controller #(parameter MASTER_CLK_FREQ = 50_000_000)
(
    // System clock and control signals
    input logic i_clk,        // System clock (typically 50MHz)
    input logic i_rst,        // Asynchronous reset (active high)
    input logic i_ena,        // Module enable (active high)
    input logic i_stb,        // Strobe signal (not used in final version)
    
    // UART interface signals for RS485 communication
    input logic i_uart_rx,    // Serial data received from JVS device
    output logic o_uart_tx,   // Serial data transmitted to JVS device
    input logic i_sense,      // JVS SENSE line (read-only for master)
    output logic o_rx485_dir, // RS485 transceiver direction control (0=RX, 1=TX)
    
    // Output registers compatible with Analogue Pocket SNAC format
    output logic [15:0] p1_btn_state,   // Player 1 button states
    output logic [31:0] p1_joy_state,   // Player 1 analog stick states
    output logic [15:0] p2_btn_state,   // Player 2 button states
    output logic [31:0] p2_joy_state,   // Player 2 analog stick states
    output logic [15:0] p3_btn_state,   // Player 3 button states (reserved)
    output logic [15:0] p4_btn_state,    // Player 4 button states (reserved)
    
    // Screen position outputs (light gun/touch screen) - raw 16-bit data
    output logic [15:0] screen_pos_x,   // Screen X position (16-bit from JVS)
    output logic [15:0] screen_pos_y,   // Screen Y position (16-bit from JVS)
    output logic has_screen_pos,        // Device supports screen position inputs

    // Coin counter outputs (up to 4 coin slots)
    output logic [15:0] coin_count[4],  // Coin counters for each slot (16-bit values)
    output logic coin1,                 // Coin increase signal for slot 1
    output logic coin2,                 // Coin increase signal for slot 2
    output logic coin3,                 // Coin increase signal for slot 3
    output logic coin4,                 // Coin increase signal for slot 4
    
    // GPIO control from SNAC
    input logic [7:0] gpio_output_value, // GPIO output value from SNAC (0x80=active, 0x00=inactive)

    //JVS node information structure
    output logic jvs_data_ready,
    output jvs_node_info_t jvs_nodes,
    //RAM interface for node names (for debug/display purposes)
    output logic [7:0] node_name_rd_data,
    input logic [6:0] node_name_rd_addr
); 

    localparam UART_CLKS_PER_BIT = MASTER_CLK_FREQ / 115200;
//==================================================================================
// Show in Quartus Synthesis if dummy data is used for simulation without JVS device
//==================================================================================
`ifdef USE_DUMMY_JVS_DATA
  initial $warning("=== USE_DUMMY_JVS_DATA is defined (=%0d). Using DUMMY data for JVS IO device ===", `USE_DUMMY_JVS_DATA);
`else
  initial $warning("=== USE_DUMMY_JVS_DATA is NOT defined.  Using REAL data for JVS IO device ===");
`endif

    //=========================================================================
    // JVS_COM INTERFACE SIGNALS (New modular interface)
    //=========================================================================
    // These signals will be used to communicate with the jvs_com module
    
    // TX interface signals
    logic [7:0] com_tx_data;        // Data byte to transmit  
    logic       com_tx_data_push;   // Pulse to push TX data
    logic       com_tx_cmd_push;    // Pulse to push TX command (stores in FIFO)
    logic [7:0] com_dst_node;       // Destination node address
    logic       com_commit;         // Pulse to commit and transmit frame
    logic       com_tx_ready;       // TX ready to accept data
    
    // RX interface signals
    logic [7:0] com_rx_byte;        // Current data byte from RX
    logic       com_rx_next;        // Pulse to get next RX byte
    logic [7:0] com_rx_remaining;   // Bytes remaining (0 = current is last)
    logic [7:0] com_src_node;       // Source node of response
    logic [7:0] com_src_cmd;        // CMD from command FIFO
    logic [7:0] com_src_cmd_status; // Status of src_cmd (STATUS_NORMAL/STATUS_BUSY)
    logic       com_src_cmd_next;   // Pulse to get next command from FIFO
    logic [4:0] com_src_cmd_count;  // Number of commands available in FIFO
    logic       com_rx_complete;    // Pulse when RX frame complete
    logic       com_rx_error;       // RX checksum or format error

    // Debug/Status signals from jvs_com
    logic [3:0] com_tx_state_debug;
    logic [3:0] com_rx_state_debug;
    logic [7:0] com_frames_tx_count;
    logic [7:0] com_frames_rx_count;
    logic [7:0] com_checksum_errors_count;

    // Edge detection for RX complete signal
    logic       com_rx_complete_d;      // Delayed version for edge detection
    wire        com_rx_complete_negedge = com_rx_complete_d & ~com_rx_complete;

    // Name copying variables for device identification parsing
    logic [7:0] copy_write_idx;         // Write index for name copying
   
    logic [3:0] current_player;
    logic [7:0] current_channel;
    //=========================================================================
    // JVS COMMUNICATION MODULE INSTANCE
    //=========================================================================
    
    // Instantiate JVS communication module
    jvs_com #(
        .MASTER_CLK_FREQ(MASTER_CLK_FREQ),
        .JVS_BUFFER_SIZE(256)
    ) jvs_com_inst (
        .clk_sys(i_clk),  // RX_NEXT/TX_NEXT states handle timing control
        .reset(i_rst),
        .i_ena(i_ena),

        // UART Physical Interface
        .uart_rx(i_uart_rx),
        .uart_tx(o_uart_tx),
        .o_rs485_dir(o_rx485_dir),          // RS485 direction control (active-high)
        
        // TX Interface
        .tx_data(com_tx_data),
        .tx_data_push(com_tx_data_push),
        .tx_cmd_push(com_tx_cmd_push),
        .dst_node(com_dst_node),
        .commit(com_commit),
        .tx_ready(com_tx_ready),
        
        // RX Interface
        .rx_byte(com_rx_byte),
        .rx_next(com_rx_next),
        .rx_remaining(com_rx_remaining),
        .src_node(com_src_node),
        .src_cmd(com_src_cmd),
        .src_cmd_status(com_src_cmd_status),
        .src_cmd_next(com_src_cmd_next),
        .src_cmd_count(com_src_cmd_count),
        .rx_complete(com_rx_complete),
        .rx_error(com_rx_error),
        
        // Debug/Status Interface (unused for now)
        .tx_state_debug(com_tx_state_debug),
        .rx_state_debug(com_rx_state_debug),
        .frames_tx_count(com_frames_tx_count),
        .frames_rx_count(com_frames_rx_count),
        .checksum_errors_count(com_checksum_errors_count)
    );
    
    // RS485 direction is now directly connected to jvs_com output

    //=========================================================================
    // JVS PROTOCOL CONSTANTS
    //=========================================================================

    // Common delay timings (in clock cycles at MASTER_CLK_FREQ)
    localparam logic [31:0] INIT_DELAY_COUNT = MASTER_CLK_FREQ * 5.4; // 5.4 seconds
    localparam logic [31:0] FIRST_RESET_DELAY_COUNT = MASTER_CLK_FREQ * 2; // 2 seconds
    localparam logic [31:0] SECOND_RESET_DELAY_COUNT = MASTER_CLK_FREQ / 2; // 0.5 seconds
    localparam logic [15:0] TX_SETUP_DELAY_COUNT = MASTER_CLK_FREQ / 100_000; // ~10µs
    localparam logic [15:0] TX_HOLD_DELAY_COUNT = MASTER_CLK_FREQ / 33_333; // ~30µs
    localparam logic [31:0] RX_TIMEOUT_COUNT = MASTER_CLK_FREQ * 2; // 1s (augmenté pour le parsing des features)
    localparam logic [31:0] POLL_INTERVAL_COUNT = MASTER_CLK_FREQ / 1_000; // 1ms
    localparam logic [31:0] SETADDR_TO_IOIDENT_DELAY = MASTER_CLK_FREQ / 500; // 2ms delay after SETADDR
    localparam logic [31:0] IOIDENT_TO_CMDREV_DELAY = MASTER_CLK_FREQ / 1000; // 1ms delay after IOIDENT
    localparam logic [31:0] CMDREV_TO_JVSREV_DELAY = MASTER_CLK_FREQ / 1000; // 1ms delay after CMDREV
    localparam logic [31:0] JVSREV_TO_COMMVER_DELAY = MASTER_CLK_FREQ / 1000; // 1ms delay after JVSREV
    localparam logic [31:0] COMMVER_TO_FEATURES_DELAY = MASTER_CLK_FREQ / 1000; // 1ms delay after COMMVER
    localparam logic [31:0] FEATURES_TO_IDLE_DELAY = MASTER_CLK_FREQ / 500; // 2ms delay after FEATURES
    localparam logic [31:0] POLLING_INTERVAL_DELAY = MASTER_CLK_FREQ / 1000; // 1ms delay between polling cycles


    //=========================================================================
    // JVS COMMAND DEFINITIONS (Based on JVS Specification)
    //=========================================================================
    
    // Standard JVS protocol bytes
    localparam JVS_SYNC_BYTE = 8'hE0;        // Frame start synchronization byte
    localparam JVS_BROADCAST_ADDR = 8'hFF;   // Broadcast address for all devices
    localparam JVS_HOST_ADDR = 8'h00;        // Host/Master address
    
    // Global Commands - Work with any device address or broadcast (0xFF)
    localparam CMD_RESET = 8'hF0;            // [F0 D9] Reset all devices on bus
                                             // Args: D9 (fixed argument)
                                             // Response: No response (devices reset)
    localparam CMD_RESET_ARG = 8'hD9;        // Argument byte that must follow CMD_RESET
    
    localparam CMD_SETADDR = 8'hF1;          // [F1 addr] Assign address to device
                                             // Args: addr (1-31, device address)
                                             // Response: [report] - report=01 if success
    
    localparam CMD_COMMCHG = 8'hF2;          // [F2 baudrate] Change communication speed
                                             // Args: baudrate (communication speed code)
                                             // Response: [report] - report=01 if success
    
    // Initialize Commands - Device identification and capability discovery
    localparam CMD_IOIDENT = 8'h10;          // [10] Read device identification string
                                             // Args: none
                                             // Response: [report name_string 00]
                                             //   name_string: ASCII device name (manufacturer;product;version;region,comment)
    
    localparam CMD_CMDREV = 8'h11;           // [11] Read command format revision
                                             // Args: none  
                                             // Response: [report revision]
                                             //   revision: BCD format (e.g. 0x13 for v1.3)
    
    localparam CMD_JVSREV = 8'h12;           // [12] Read JVS specification revision
                                             // Args: none
                                             // Response: [report revision]
                                             //   revision: BCD format (e.g. 0x30 for v3.0)
    
    localparam CMD_COMMVER = 8'h13;          // [13] Read communication version
                                             // Args: none
                                             // Response: [report version]
                                             //   version: BCD format (e.g. 0x10 for v1.0)
    
    localparam CMD_FEATCHK = 8'h14;          // [14] Check device features/capabilities
                                             // Args: none
                                             // Response: [report func_data... 00]
                                             //   func_data: loop of 4-byte blocks [func_code param1 param2 param3] loop end with 00
    
    localparam CMD_MAINID = 8'h15;           // [15] Send main board ID to I/O device
                                             // Args: [main_pcb_id_string 00] - ASCII string up to 100 chars
                                             //   Format: "Maker;Game;Version;Details" separated by semicolons
                                             //   Example: "NAMCO LTD.;TEKKEN2;ver1.6; TEKKEN2 ver B"
                                             // Response: [report] - report=01 if success
    
    // Data I/O Commands - Input reading and data retrieval
    localparam CMD_SWINP = 8'h20;            // [20 players bytes] Read switch inputs (digital buttons)
                                             // Args: players (number of players), bytes (total bytes needed for bits per player)
                                             // Response: [report switch_data...]
                                             //   switch_data: players × bytes of digital input data
    
    localparam CMD_COININP = 8'h21;          // [21 slots] Read coin inputs and counter
                                             // Args: slots (number of coin slots to read)
                                             // Response: [report coin_status...]
                                             //   coin_status: loop of 2 bytes [condition(2 bits) counter_MSB(6 bits) counter_LSB]
    
    // Coin Input Condition Codes (Table 12)
    localparam COIN_CONDITION_NORMAL = 2'b00;        // Normal operation
    localparam COIN_CONDITION_JAM = 2'b01;           // Coin jam detected
    localparam COIN_CONDITION_DISCONNECTED = 2'b10;  // Coin mechanism disconnected  
    localparam COIN_CONDITION_BUSY = 2'b11;          // Coin mechanism busy

    localparam CMD_ANLINP = 8'h22;           // [22 channels] Read analog inputs
                                             // Args: channels (number of analog channels)
                                             // Response: [report analog_data...]
                                             //   analog_data: 2 bytes per channel [data_MSB data_LSB]
    
    localparam CMD_ROTINP = 8'h23;           // [23 channels] Read rotary inputs
                                             // Args: channels (number of rotary channels to read)
                                             // Response: [report rotary_data...]
                                             //   rotary_data: 2 bytes per channel [data_MSB data_LSB]
    
    localparam CMD_KEYINP = 8'h24;           // [24] Read keycode inputs
                                             // Args: none
                                             // Response: [report keycode]
                                             //   keycode: ASCII key code or 00 if no key
    
    localparam CMD_SCRPOSINP = 8'h25;        // [25 channels] Read screen position inputs (light gun/touch)
                                             // Args: channel index to read
                                             // Response: [report pos_data...]
                                             //   pos_data: 4 bytes [x_MSB x_LSB y_MSB y_LSB]
    
    localparam CMD_MISCSWINP = 8'h26;        // [26 bytes] Read miscellaneous switch inputs
                                             // Args: bytes (number of misc input bytes, depends on bits defined in feature check)
                                             // Response: [report misc_data...]
                                             //   misc_data: specified number of misc input bytes

    localparam CMD_PAYCNT = 8'h2E;           // [2E channel_index] Payout coins/tokens aka. redemption
                                             // Args: channel_index
                                             // Response: [report hopper_status remaining_hi remaining_mid remaining_low]

    localparam CMD_RETRANSMIT = 8'h2F;       // [2F] Retransmit previous response
                                             // Args: none
                                             // Response: Previous response is retransmitted

    localparam CMD_COINDEC = 8'h30;          // [30 slots_index amount_msb amount_lsb] Decrease selected coin counter of specified value
                                             // Args: slot_index, amount_msb, amount_lsb
                                             // Response: [report] - report=01 if success

    localparam CMD_PAYINC = 8'h31;           // [31 slots payval...] Increase payout counters
                                             // Args: slots (number of payout slots), payval per slot (increase amount)
                                             // Response: [report] - report=01 if success
    
    localparam CMD_OUTPUT1 = 8'h32;          // [32 bytes data...] General purpose output 1
                                             // Args: bytes (number of output bytes), data per byte
                                             // Response: [report] - report=01 if success
    
    localparam CMD_ANLOUT = 8'h33;           // [33 channels data...] Analog output control
                                             // Args: channels (number of analog outputs), 2 bytes data per channel [MSB LSB]
                                             // Response: [report] - report=01 if success
    
    localparam CMD_CHAROUT = 8'h34;          // [34 line pos string...] Character display output
                                             // Args: line (display line), pos (position), string data
                                             // Response: [report] - report=01 if success
    
    localparam CMD_COININC = 8'h35;          // [35 slots incval...] Increase coin counters
                                             // Args: slots (number of coin slots), incval per slot (increase amount)
                                             // Response: [report] - report=01 if success
    
    localparam CMD_PAYDEC = 8'h36;           // [36 slots decval...] Decrease payout counters
                                             // Args: slots (number of payout slots), decval per slot (decrease amount)
                                             // Response: [report] - report=01 if success
    
    localparam CMD_OUTPUT2 = 8'h37;          // [37 bytes data...] General purpose output 2
                                             // Args: bytes (number of output bytes), data per byte
                                             // Response: [report] - report=01 if success
    
    localparam CMD_OUTPUT3 = 8'h38;          // [38 bytes data...] General purpose output 3
                                             // Args: bytes (number of output bytes), data per byte
                                             // Response: [report] - report=01 if success
    

    // Status Codes - General response status (position 3 in frame)
    localparam STATUS_NORMAL = 8'h01;        // Normal operation status
    localparam STATUS_UNKNOWN_CMD = 8'h02;   // Unknown command received  
    localparam STATUS_SUM_ERROR = 8'h03;     // Checksum error in received data
    localparam STATUS_ACK_OVERFLOW = 8'h04;  // Acknowledgment overflow
    localparam STATUS_BUSY = 8'h05;          // Device busy, cannot process command
    
    // Report Codes - Command-specific status (position 4+ in frame)
    localparam REPORT_NORMAL = 8'h01;        // Normal operation
    localparam REPORT_PARAM_ERROR_COUNT = 8'h02; // Parameter error (incorrect number)
    localparam REPORT_PARAM_ERROR_DATA = 8'h03;  // Parameter error (invalid data)
    localparam REPORT_BUSY = 8'h04;          // Busy (cannot receive more commands)  

    // JVS Escape sequence constants for data byte escaping
    localparam JVS_ESCAPE_BYTE = 8'hD0;      // Escape marker byte
    localparam JVS_ESCAPED_E0 = 8'hDF;       // E0 becomes D0 DF
    localparam JVS_ESCAPED_D0 = 8'hCF;       // D0 becomes D0 CF
    
    // Function Codes - Used in feature check responses
    localparam FUNC_INPUT_DIGITAL = 8'h01;    // [01 players bytesperplayer unused] Digital inputs
    localparam FUNC_INPUT_COIN = 8'h02;       // [02 slots unused unused] Coin inputs
    localparam FUNC_INPUT_ANALOG = 8'h03;     // [03 channels bits unused] Analog inputs (channels×bits resolution)
    localparam FUNC_INPUT_ROTARY = 8'h04;     // [04 channels unused unused] Rotary encoder inputs
    localparam FUNC_INPUT_KEYCODE = 8'h05;    // [05 unused unused unused] Keycode inputs
    localparam FUNC_INPUT_SCREEN_POS = 8'h06; // [06 channels bits unused] Screen position inputs (channels×bits)
    localparam FUNC_INPUT_MISC_DIGITAL = 8'h07; // [07 bytes unused unused] Miscellaneous digital inputs
    localparam FUNC_OUTPUT_CARD = 8'h10;      // [10 slots unused unused] Card system outputs
    localparam FUNC_OUTPUT_HOPPER = 8'h11;    // [11 slots unused unused] Medal/token hopper outputs  
    localparam FUNC_OUTPUT_DIGITAL = 8'h12;   // [12 bytes unused unused] Digital outputs (lights/solenoids)
    localparam FUNC_OUTPUT_ANALOG = 8'h13;    // [13 channels unused unused] Analog outputs
    localparam FUNC_OUTPUT_CHAR = 8'h14;      // [14 lines columns type] Character display outputs
    localparam FUNC_OUTPUT_BACKUP = 8'h15;    // [15 unused unused unused] Backup data support

    localparam JVS_FUNC_LENGTH = 8'd4;          // Each function block is 4 bytes long
    
    // Character Output Type codes (Table 9)
    localparam JVS_CHAR_TYPE_UNKNOWN = 8'h00;           // Unknown
    localparam JVS_CHAR_TYPE_ASCII_NUMERIC = 8'h01;     // ASCII (numeric)
    localparam JVS_CHAR_TYPE_ASCII_ALPHANUM = 8'h02;    // ASCII (alphanumeric)
    localparam JVS_CHAR_TYPE_ASCII_KATAKANA = 8'h03;    // ASCII (alphanumeric, half-width katakana)
    localparam JVS_CHAR_TYPE_ASCII_KANJI = 8'h04;       // ASCII (kanji support, SHIFT-JIS)
    
    // JVS Frame structure constants for better code readability
    localparam JVS_SYNC_POS = 8'd0;          // Position of sync byte (E0)
    localparam JVS_ADDR_POS = 8'd1;          // Position of address byte
    localparam JVS_LENGTH_POS = 8'd2;        // Position of length byte
    localparam JVS_DATA_START = 8'd4;        // Start position of data bytes (RX) - after status and include report bytes
    localparam JVS_STATUS_POS = 8'd3;        // Position of status byte in response
    localparam JVS_REPORT_POS = 8'd4;        // Position of report byte in response (should be processed)
    localparam JVS_CMD_START = 8'd3;         // Start position of command bytes (TX)
    localparam JVS_OVERHEAD = 8'd2;          // Overhead for length calculation (includes checksum + command byte)
    localparam JVS_CHECKSUM_SIZE = 8'd1;     // Checksum is coded on one byte

    // Buffer size configuration for resource optimization
    localparam RX_BUFFER_SIZE = 128;         // Size of RX buffers (I/O Identify max 106 bytes)
    localparam TX_BUFFER_SIZE = 24;          // Size of TX buffer (max frame ~21 bytes)
    
    // JVS node management constants
    //localparam MAX_JVS_NODES = 2;            // Maximum supported JVS nodes (current implementation)
    //localparam NODE_NAME_SIZE = 100;         // Maximum size for node identification strings (per JVS spec)
    // Defined in jvs_node_info_pkg.sv

    //=========================================================================
    // STATE MACHINE DEFINITIONS
    //=========================================================================
    
    //=========================================================================
    // MAIN JVS PROTOCOL STATE MACHINE (6-bit states)
    // Controls overall JVS protocol sequence from initialization to input polling
    //=========================================================================
    
    // INITIALIZATION SEQUENCE STATES (5.4s + 2s + 0.5s delays)
    localparam STATE_IDLE = 6'h00;             // Idle state - continuous input polling (1ms interval)
    localparam STATE_INIT_DELAY = 6'h02;       // Initial 5.4s delay for system stabilization
    localparam STATE_FIRST_RESET = 6'h03;      // Send first reset command (F0 D9)
    localparam STATE_FIRST_RESET_DELAY = 6'h04; // 2-second delay after first reset
    localparam STATE_SECOND_RESET = 6'h05;     // Send second reset command for reliability
    localparam STATE_SECOND_RESET_DELAY = 6'h06; // 0.5-second delay after second reset
    
    // DEVICE DISCOVERY SEQUENCE STATES
    localparam STATE_SEND_SETADDR = 6'h07;     // Send address assignment command (F1 01)
    localparam RX_PARSE_SETADDR = 6'h08;    // Parse address assignment response
    localparam STATE_SEND_IOIDENT = 6'h09;     // Send device identification request (10)
    localparam RX_PARSE_IOIDENT = 6'h0A;    // Parse device ID string response
    localparam STATE_SEND_CMDREV = 6'h0B;      // Send command revision request (11)
    localparam RX_PARSE_CMDREV = 6'h0C;     // Parse command revision response (BCD format)
    localparam STATE_SEND_JVSREV = 6'h0D;      // Send JVS revision request (12)
    localparam RX_PARSE_COMMVER = 6'h0E;    // Parse communications version response (BCD format)
    localparam RX_PARSE_JVSREV = 6'h0F;     // Parse JVS revision response (BCD format)
    localparam STATE_SEND_COMMVER = 6'h10;     // Send communications version request (13)
    localparam STATE_SEND_FEATCHK = 6'h11;     // Send feature check request (14)
    
    // GENERIC FLOW CONTROL STATES
    localparam STATE_WAIT_RX = 6'h01;          // Wait for device response with 1s timeout
    localparam STATE_MAIN_TIMER_DELAY = 6'h3D; // Generic timer delay state - returns to return_state when done
    
    // INPUT POLLING SEQUENCE STATES (chained command construction)
    localparam STATE_SEND_INPUTS = 6'h12;         // Start input polling sequence
    localparam STATE_SEND_INPUTS_SWITCH = 6'h13;  // Add switch/button inputs (20) if available
    localparam STATE_SEND_INPUTS_COIN = 6'h14;    // Add coin inputs (21) if available
    localparam STATE_SEND_INPUTS_ANALOG = 6'h15;  // Add analog inputs (22) if available (joysticks)
    localparam STATE_SEND_INPUTS_ROTARY = 6'h16;  // Add rotary inputs (23) if available
    localparam STATE_SEND_INPUTS_KEYCODE = 6'h17; // Add keycode inputs (24) if available
    localparam STATE_SEND_INPUTS_SCREEN = 6'h18;  // Add screen position (25) if available (light gun)
    localparam STATE_SEND_INPUTS_MISC = 6'h19;    // Add misc inputs (26) if available
    localparam STATE_SEND_OUTPUT_DIGITAL = 6'h1A; // Send digital output command (32) for GPIO
    localparam STATE_SEND_OUTPUT_ANALOG = 6'h3E; // Send analog output command (33) for GPIO
    localparam STATE_SEND_FINALIZE = 6'h1B;       // Finalize chained command frame and transmit
    
    // RESET ARGUMENT STATES (for double reset sequence)
    localparam STATE_FIRST_RESET_ARG = 6'h1C;     // Push first reset argument (D9) and commit
    localparam STATE_SECOND_RESET_ARG = 6'h1D;    // Push second reset argument (D9) and commit
    
    // GENERIC HELPER STATES
    localparam STATE_TX_NEXT = 6'h1E;             // Generic TX byte advance state
    localparam STATE_RX_NEXT = 6'h1F;             // Generic RX byte advance state
    localparam STATE_FATAL_ERROR = 6'h20;         // Fatal error state - stops execution

    //=========================================================================
    // RX PARSING STATES (6-bit states for complex response handling)
    // These states handle parsing of JVS command responses
    //=========================================================================
    
    // FEATURE PARSING STATES
    localparam RX_PARSE_FEATURES = 6'h21;      // Parse device feature/capability data (14 response)
    localparam RX_PARSE_FEATURES_FUNCS = 6'h22; // Parse individual function capabilities
    localparam RX_PARSE_FUNC_DIGITAL = 6'h23;  // Parse digital input function parameters
    localparam RX_PARSE_FUNC_COIN = 6'h24;     // Parse coin input function parameters
    localparam RX_PARSE_FUNC_ANALOG = 6'h25;   // Parse analog input function parameters
    localparam RX_PARSE_FUNC_ROTARY = 6'h26;   // Parse rotary input function parameters
    localparam RX_PARSE_FUNC_SCREEN = 6'h27;   // Parse screen position function parameters
    localparam RX_PARSE_FUNC_MISC = 6'h28;     // Parse misc digital function parameters

    localparam RX_PARSE_FUNC_CARD = 6'h29;         // Parse card system function parameters
    localparam RX_PARSE_FUNC_HOPPER = 6'h2A;       // Parse hopper function parameters
    localparam RX_PARSE_FUNC_OUT_DIGITAL = 6'h2B;  // Parse output digital function parameters
    localparam RX_PARSE_FUNC_OUT_ANALOG = 6'h2C;   // Parse output analog function parameters
    localparam RX_PARSE_FUNC_CHAR = 6'h2D;         // Parse character display function parameters

    // INPUT DATA PARSING STATES (chained command response handling)
    localparam RX_PARSE_INPUTS_START = 6'h30;   // Initialize chained input response parsing
    localparam RX_PARSE_INPUT_CMD = 6'h31;      // Dispatch to parser based on command in FIFO
    localparam RX_PARSE_INPUTS_COMPLETE = 6'h3C; // Complete chained parsing, return to polling

    // DATA I/O COMMANDS
    localparam RX_PARSE_SWINP = 6'h32;          // Parse switch/button inputs (20) response
    localparam RX_PARSE_SWINP_PLAYER = 6'h33;   // Parse per-player switch data (recursive)
    localparam RX_PARSE_COININP = 6'h34;        // Parse coin inputs (21) response
    localparam RX_PARSE_ANLINP = 6'h35;         // Parse analog inputs (22) response
    localparam RX_PARSE_ANLINP_DATA = 6'h36;    // Parse per-channel analog data (recursive)
    localparam RX_PARSE_ROTINP = 6'h37;         // Parse rotary inputs (23) response
    localparam RX_PARSE_KEYINP = 6'h38;         // Parse keycode inputs (24) response
    localparam RX_PARSE_SCRPOSINP = 6'h39;      // Parse screen position (25) response (light gun)
    localparam RX_PARSE_MISCSWINP = 6'h3A;      // Parse misc digital inputs (26) response
    // OUTPUT COMMANDS
    localparam RX_PARSE_OUTPUT1 = 6'h3B;        // Parse digital output (32) response
    
    
    
    //=========================================================================
    // STATE VARIABLES AND CONTROL REGISTERS
    //=========================================================================
    // Current state for main protocol state machine
    logic [5:0] main_state;        // Main protocol state (6-bit for extended states)
    
    // TX state management for sequential byte transmission
    logic [5:0] return_state;      // State to return to after TX_NEXT (6-bit for extended states)
    logic [7:0] cmd_pos;           // Position in current command sequence (was [2:0] - caused overflow)
    logic [3:0] current_coin;      // Current coin slot being parsed (0-3)
    
    // Temporary variables for coin parsing
    logic [1:0] temp_coin_condition;
    logic [5:0] temp_counter_msb;
    
    // Timing and protocol control
    logic [31:0] delay_counter;    // Multi-purpose delay counter
    logic [31:0] timeout_counter;  // Timeout counter for waiting states
    logic [31:0] poll_timer;       // Timer for input polling frequency
    logic [7:0] current_device_addr; // Address assigned to JVS device (usually 0x01)

    // Feature parsing control
    logic [7:0] current_func_code; // Store current function being parsed  
    
    //=========================================================================
    // JVS NODE INFORMATION STRUCTURES
    //=========================================================================
    // Structure to store information about each JVS node
    jvs_node_info_t jvs_nodes_r;

//see comments in JVS_Debugger.qsf under [JVS project settings] 
`ifdef USE_DUMMY_JVS_DATA
	jvs_node_info_t jvs_nodes_r2;
	 
    localparam jvs_node_info_t JVS_INFO_INIT = '{
        node_id: '{8'h01, 8'h02},
        node_cmd_ver: '{8'h13, 8'h11}, 
        node_jvs_ver: '{8'h30, 8'h30},  
        node_com_ver: '{8'h10, 8'h10},
        // Initialize dummy capabilities based on typical JVS device
        node_players: '{4'h2, 4'h1},              // 2 players for first device, 1 for second
        node_buttons: '{8'h0D, 8'h06},            // 13 buttons for P1, 6 for P2
        node_analog_channels: '{4'h2, 4'h0},      // 2 analog channels for first device
        node_analog_bits: '{8'h0A, 8'h08},        // 10-bit analog for first device, 8-bit for second
        node_rotary_channels: '{4'h0, 4'h0},      // No rotary encoders
        node_coin_slots: '{4'h2, 4'h1},           // 2 coin slots for first device, 1 for second
        // Additional input capabilities
        node_has_keycode_input: '{1'b0, 1'b0},    // No keycode input
        node_has_screen_pos: '{1'b0, 1'b0},       // No screen position input
        node_screen_pos_x_bits: '{8'h00, 8'h00},  // No screen X resolution
        node_screen_pos_y_bits: '{8'h00, 8'h00},  // No screen Y resolution  
        node_misc_digital_inputs: '{16'h0000, 16'h0000}, // No misc digital inputs (16-bit)
        // Output capabilities
        node_digital_outputs: '{8'h08, 8'h00},    // 8 digital outputs for first device
        node_analog_output_channels: '{4'h2, 4'h0}, // 2 analog output channels for first device
        node_card_system_slots: '{8'h00, 8'h00},  // No card system slots
        node_medal_hopper_channels: '{8'h00, 8'h00}, // No medal hopper channels
        node_has_char_display: '{1'b0, 1'b0},     // No character display
        node_char_display_width: '{8'h00, 8'h00}, // No character display width
        node_char_display_height: '{8'h00, 8'h00}, // No character display height
        node_char_display_type: '{8'h00, 8'h00},   // No character display type
        node_has_backup: '{1'b0, 1'b0}            // No backup support
    };
    assign jvs_nodes = jvs_nodes_r2;
`else 
    assign jvs_nodes = jvs_nodes_r;
`endif

    //=========================================================================
    // RAM for current node name during reception
    (* ramstyle = "M10K" *) logic [7:0] node_name_ram [0:jvs_node_info_pkg::NODE_NAME_SIZE -1];

////initial content for simulation without JVS device
`ifdef USE_DUMMY_JVS_DATA
    initial begin
        $readmemh("jvs_device_name.mem", node_name_ram); //null terminated string "namco ltd.;NAJV2;Ver1.00;JPN,Multipurpose."
    end
`endif

    //infer simple dual-port RAM for node name reading
    always_ff @(posedge i_clk) begin
        node_name_rd_data <= node_name_ram[node_name_rd_addr];
    end

    //=========================================================================
    // JVS DATA READY SIGNAL
    //=========================================================================
    logic jvs_data_ready_init, jvs_data_ready_joy;
    assign jvs_data_ready = jvs_data_ready_init | jvs_data_ready_joy;
    
    //=========================================================================
    // MAIN STATE MACHINE - JVS PROTOCOL HANDLER
    //=========================================================================
    // Implements the complete JVS initialization sequence and input polling
    
    always @(posedge i_clk) begin

        jvs_data_ready_init <= 1'b0;

        // Update delayed register for edge detection
        com_rx_complete_d <= com_rx_complete;

        // Default: Clear all jvs_com control signals (they are pulses)
        com_tx_data_push <= 1'b0;
        com_tx_cmd_push <= 1'b0;
        com_commit <= 1'b0;
        com_rx_next <= 1'b0;
        com_src_cmd_next <= 1'b0;

        if (i_rst || !i_ena) begin
            // Initialize all state variables on reset
            main_state <= STATE_INIT_DELAY;
            delay_counter <= 32'h0;
            timeout_counter <= 32'h0;
            poll_timer <= 32'h0;
            current_device_addr <= 8'h01;    // Standard JVS device address
            
            // Initialize TX state management
            return_state <= 6'h0;
            cmd_pos <= 8'h0;
            
            // Initialize jvs_com control signals
            com_tx_data <= 8'h00;
            com_tx_data_push <= 1'b0;
            com_tx_cmd_push <= 1'b0;
            com_dst_node <= 8'h00;
            com_commit <= 1'b0;
            com_rx_next <= 1'b0;
            com_src_cmd_next <= 1'b0;

            // Initialize output button and joystick states
            p1_btn_state <= 16'h0000;           // All buttons released
            p1_joy_state <= 32'h80808080;       // Analog sticks centered (0x80 = center)
            p2_btn_state <= 16'h0000;
            p2_joy_state <= 32'h80808080;
            p3_btn_state <= 16'h0000;
            p4_btn_state <= 16'h0000;

            // Initialize coin counters
            coin_count[0] <= 16'h0000;
            coin_count[1] <= 16'h0000;
            coin_count[2] <= 16'h0000;
            coin_count[3] <= 16'h0000;

            // Initialize JVS node information (single node only)
            jvs_nodes_r.node_id[0] <= 8'h01;
            jvs_nodes_r.node_cmd_ver[0] <= 8'h00;
            jvs_nodes_r.node_jvs_ver[0] <= 8'h00;
            jvs_nodes_r.node_com_ver[0] <= 8'h00;
            jvs_nodes_r.node_players[0] <= 4'h0;
            jvs_nodes_r.node_buttons[0] <= 8'h0;
            jvs_nodes_r.node_analog_channels[0] <= 4'h0;
            jvs_nodes_r.node_rotary_channels[0] <= 4'h0;
            // Additional input capabilities (not yet supported)
            jvs_nodes_r.node_has_keycode_input[0] <= 1'b0;
            jvs_nodes_r.node_has_screen_pos[0] <= 1'b0;
            jvs_nodes_r.node_screen_pos_x_bits[0] <= 8'h0;
            jvs_nodes_r.node_screen_pos_y_bits[0] <= 8'h0;
            // Initialize has_screen_pos output
            has_screen_pos <= 1'b0;
            jvs_nodes_r.node_misc_digital_inputs[0] <= 16'h0;
            // Output capabilities
            jvs_nodes_r.node_digital_outputs[0] <= 8'h0;
            jvs_nodes_r.node_analog_output_channels[0] <= 4'h0;
            jvs_nodes_r.node_card_system_slots[0] <= 8'h0;
            jvs_nodes_r.node_medal_hopper_channels[0] <= 8'h0;
            jvs_nodes_r.node_has_char_display[0] <= 1'b0;
            jvs_nodes_r.node_char_display_width[0] <= 8'h0;
            jvs_nodes_r.node_char_display_height[0] <= 8'h0;
            jvs_nodes_r.node_char_display_type[0] <= 8'h0;
            jvs_nodes_r.node_has_backup[0] <= 1'b0;

            // Initialize edge detection register
            com_rx_complete_d <= 1'b0;
        end else begin
            case (main_state)
                //-------------------------------------------------------------
                // IDLE STATE - Continuous input polling for responsive gaming
                //-------------------------------------------------------------
                STATE_IDLE: begin
                    
                    // Fast polling timer for inputs - 1ms interval
                    // This provides responsive gaming experience with minimal latency
                    //if (poll_timer < 32'h0C350) begin  // 50,000 cycles = 1ms at 50MHz
                    if (poll_timer < POLL_INTERVAL_COUNT) begin  // 1ms
                        poll_timer <= poll_timer + 1;
                    end else begin
                        poll_timer <= 32'h0;
                        main_state <= STATE_SEND_INPUTS;
                    end
                end

                //-------------------------------------------------------------
                // INITIALIZATION DELAY - Wait for system stabilization
                //-------------------------------------------------------------
                STATE_INIT_DELAY: begin
                    // Initial delay for core I/O initialization - 5.4 seconds
                    // This ensures the FPGA core and external circuits are fully stable
                    //if (delay_counter < 32'h10000000) begin  // 268,435,456 cycles ≈ 5.4s at 50MHz
                    if (delay_counter < INIT_DELAY_COUNT) begin  // 5.4 seconds
                        delay_counter <= delay_counter + 1;
                    end else begin
                        delay_counter <= 32'h0;
                        main_state <= STATE_FIRST_RESET;
                    end
                end

                //-------------------------------------------------------------
                // FIRST RESET COMMAND - Begin JVS device initialization
                //-------------------------------------------------------------
                STATE_FIRST_RESET: begin
                    // Send first RESET command using sequential byte transmission
                    // JVS requires two reset commands for reliable initialization
                    if (com_tx_ready) begin
                        com_dst_node <= JVS_BROADCAST_ADDR;  // FF - Broadcast to all devices
                        return_state <= STATE_FIRST_RESET;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_RESET;     // Reset command (0xF0)
                                com_tx_data_push <= 1'b1;     // Push as data because RESET does not give answer
                                main_state <= STATE_TX_NEXT; // Go to TX_NEXT
                            end
                            3'd1: begin
                                com_tx_data <= CMD_RESET_ARG; // Reset argument (0xD9)
                                com_tx_data_push <= 1'b1;    // Push as data  
                                main_state <= STATE_TX_NEXT; // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                cmd_pos <= 8'd0;
                                main_state <= STATE_FIRST_RESET_DELAY;
                            end
                        endcase
                    end
                end

                //-------------------------------------------------------------
                // DELAY AFTER FIRST RESET
                //-------------------------------------------------------------
                STATE_FIRST_RESET_DELAY: begin

                    // 2 second delay after first RESET
                    // Allows JVS devices to complete their reset sequence
                    //if (delay_counter < 32'h6000000) begin  // 100,663,296 cycles = 2s at 50MHz
                    if (delay_counter <FIRST_RESET_DELAY_COUNT) begin  //   2 seconds
                        delay_counter <= delay_counter + 1;
                    end else begin
                        delay_counter <= 32'h0;
                        main_state <= STATE_SECOND_RESET;
                    end
                end

                //-------------------------------------------------------------
                // SECOND RESET COMMAND - Ensure complete device reset
                //-------------------------------------------------------------
                STATE_SECOND_RESET: begin
                    // Send second RESET command using sequential byte transmission (identical to first)
                    if (com_tx_ready) begin
                        com_dst_node <= JVS_BROADCAST_ADDR;  // FF - Broadcast to all devices
                        return_state <= STATE_SECOND_RESET;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_RESET;     // Reset command (0xF0)
                                com_tx_data_push <= 1'b1;     // Push as data does not give answer !!
                                main_state <= STATE_TX_NEXT; // Go to TX_NEXT
                            end
                            3'd1: begin
                                com_tx_data <= CMD_RESET_ARG; // Reset argument (0xD9)
                                com_tx_data_push <= 1'b1;    // Push as data  
                                main_state <= STATE_TX_NEXT; // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                cmd_pos <= 8'd0;
                                main_state <= STATE_SECOND_RESET_DELAY;
                            end
                        endcase
                    end
                end

                //-------------------------------------------------------------
                // DELAY AFTER SECOND RESET
                //-------------------------------------------------------------
                STATE_SECOND_RESET_DELAY: begin
                    // 500ms delay after second RESET
                    // Shorter delay as devices should be ready after two resets
                    //if (delay_counter < 32'h1800000) begin  // 25,165,824 cycles = 500ms at 50MHz
                    if (delay_counter < SECOND_RESET_DELAY_COUNT) begin  // 500ms
                        delay_counter <= delay_counter + 1;
                    end else begin
                        delay_counter <= 32'h0;
                        main_state <= STATE_SEND_SETADDR;
                    end
                end

                //-------------------------------------------------------------
                // SET ADDRESS COMMAND - Assign unique address to device
                //-------------------------------------------------------------
                STATE_SEND_SETADDR: begin
                    // Send SET ADDRESS command using sequential byte transmission
                    // This assigns a unique address (0x01) to the JVS device
                    if (com_tx_ready) begin
                        $display("[CONTROLLER][STATE_SEND_SETADDR] cmd_pos 0x%02X", cmd_pos);
                        // Initialize command parameters on first entry
                        com_dst_node <= JVS_BROADCAST_ADDR;  // FF - Still broadcast for address assignment
                        return_state <= STATE_SEND_SETADDR;
                        main_state <= STATE_TX_NEXT;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_SETADDR;         // Set address command (0xF1)
                                com_tx_cmd_push <= 1'b1;            // Push as command
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            3'd1: begin
                                com_tx_data <= current_device_addr; // 01 - Address to assign
                                com_tx_data_push <= 1'b1;           // Push as data
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end
                end
                
                //-------------------------------------------------------------
                // PARSE SETADDR RESPONSE - Verify address assignment
                //-------------------------------------------------------------
                RX_PARSE_SETADDR: begin
                    $display("[CONTROLLER][RX_PARSE_SETADDR] cmd_pos 0x%02X, rx_byte 0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_SETADDR;
                    case (cmd_pos)
                        3'd0: begin
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            // Check REPORT byte
                            if (com_rx_byte == REPORT_NORMAL) begin
                                $display("[CONTROLLER][RX_PARSE_SETADDR] Address %d accepted %d", current_device_addr, com_rx_remaining);
                                com_rx_next <= 1'b1;     // Advance to first name character
                                main_state <= STATE_RX_NEXT;
                            end else begin
                                $display("[CONTROLLER][RX_PARSE_SETADDR] ERROR: Bad REPORT 0x%02X for SETADDR", com_rx_byte);
                                $display("[CONTROLLER][FATAL_ERROR] SETADDR failed - device rejected address assignment");
                                main_state <= STATE_FATAL_ERROR;
                            end
                        end
                        default: begin
                            cmd_pos <= 8'd0;          // Reset position for next command
                            // Add delay before sending IOIDENT command
                            delay_counter <= SETADDR_TO_IOIDENT_DELAY;
                            return_state <= STATE_SEND_IOIDENT;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                            $display("[CONTROLLER] SETADDR complete, adding %0d cycle delay before IOIDENT", SETADDR_TO_IOIDENT_DELAY);
                        end
                    endcase
                end
                
                //-------------------------------------------------------------
                // READ ID COMMAND - Request device identification
                //-------------------------------------------------------------
                STATE_SEND_IOIDENT: begin
                    if (com_tx_ready) begin
                        $display("[CONTROLLER][STATE_SEND_IOIDENT] cmd_pos 0x%02X", cmd_pos);
                        // Initialize command parameters on first entry
                        com_dst_node <= current_device_addr; // 01 - Address specific device
                        return_state <= STATE_SEND_IOIDENT;
                        main_state <= STATE_TX_NEXT;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_IOIDENT;          // IO identity command (0x10)
                                com_tx_cmd_push <= 1'b1;             // Push as command
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition then wait answer
                                com_commit <= 1'b1;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end
                end
                
                //-------------------------------------------------------------
                // PARSE IOIDENT RESPONSE - Extract device name
                //-------------------------------------------------------------
                RX_PARSE_IOIDENT: begin
                    return_state <= RX_PARSE_IOIDENT;
                    case (cmd_pos)
                        3'd0: begin
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            // Check REPORT byte
                            if (com_rx_byte == REPORT_NORMAL) begin
                                copy_write_idx <= 8'd0;  // Reset write index for name copying
                                com_rx_next <= 1'b1;     // Advance to first name character
                                main_state <= STATE_RX_NEXT;
                            end else begin
                                $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for IOIDENT", com_rx_byte);
                                $display("[CONTROLLER][FATAL_ERROR] IOIDENT failed - device cannot provide identification");
                                main_state <= STATE_FATAL_ERROR;
                            end
                        end
                        default: begin
                            // Copy device name characters until null terminator or end of data
                            if (com_rx_remaining > 0) begin // > 1 because we need to leave room for checksum
                                if (com_rx_byte == 8'h00) begin
                                    // Found null terminator, store it and finish copying
                                    jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= 8'h00;
                                    /*
                                    $display("[CONTROLLER][RX_PARSE_IOIDENT] Name copy complete, %d chars %d", copy_write_idx, com_rx_remaining);
                                    $write("[CONTROLLER][RX_PARSE_IOIDENT] Device name: ");
                                    for (int i = 0; i < copy_write_idx; i++) begin
                                        $write("%c", jvs_nodes_r.node_name[current_device_addr - 1][i]);
                                    end
                                    $display("");
                                    */
                                    cmd_pos <= 8'd0;  // Reset position for next command
                                    // Add delay before sending CMDREV command
                                    delay_counter <= IOIDENT_TO_CMDREV_DELAY;
                                    return_state <= STATE_SEND_CMDREV;
                                    main_state <= STATE_MAIN_TIMER_DELAY;
                                    $display("[CONTROLLER] IOIDENT complete, adding %0d cycle delay before CMDREV", IOIDENT_TO_CMDREV_DELAY);
                                end else if (copy_write_idx < jvs_node_info_pkg::NODE_NAME_SIZE - 1) begin
                                    // Copy character to node name buffer
                                    jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= com_rx_byte;
                                    copy_write_idx <= copy_write_idx + 1;
                                    com_rx_next <= 1'b1;     // Advance to first name character
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    // Buffer full, skip remaining characters until null terminator
                                    $display("[CONTROLLER][RX_PARSE_IOIDENT] Name buffer full, skipping chars");
                                    com_rx_next <= 1'b1;     // Advance to first name character
                                    cmd_pos <= 8'd0;  // Reset position for next command
                                    delay_counter <= IOIDENT_TO_CMDREV_DELAY;
                                    return_state <= STATE_SEND_CMDREV;
                                    main_state <= STATE_MAIN_TIMER_DELAY;
                                end
                            end else begin
                                // End of data reached without null terminator
                                $display("[CONTROLLER][RX_PARSE_IOIDENT] End of data reached, name copy complete");
                                cmd_pos <= 8'd0;
                                delay_counter <= IOIDENT_TO_CMDREV_DELAY;
                                return_state <= STATE_SEND_CMDREV;
                                main_state <= STATE_MAIN_TIMER_DELAY;
                            end
                        end
                    endcase
                end
                
                //-------------------------------------------------------------
                // COMMAND REVISION REQUEST - Get command format revision
                //-------------------------------------------------------------
                STATE_SEND_CMDREV: begin
                    $display("[CONTROLLER] STATE_SEND_CMDREV: com_tx_ready=%b, cmd_pos=%d", com_tx_ready, cmd_pos);
                    if (com_tx_ready) begin
                        $display("[CONTROLLER][STATE_SEND_CMDREV] cmd_pos 0x%02X", cmd_pos);
                        // Initialize command parameters on first entry
                        main_state <= STATE_TX_NEXT;
                        com_dst_node <= current_device_addr; // 01 - Address specific device
                        return_state <= STATE_SEND_CMDREV;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                $display("[CONTROLLER] Pushing CMDREV command: data=0x%02X", CMD_CMDREV);
                                com_tx_data <= CMD_CMDREV;          // Command revision command (0x11)
                                com_tx_cmd_push <= 1'b1;            // Push as command (ONLY this one!)
                                $display("[CONTROLLER] com_tx_cmd_push set to 1");
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end else begin
                        $display("[CONTROLLER] Waiting for com_tx_ready...");
                    end
                end
                
                //-------------------------------------------------------------
                // PARSE CMDREV RESPONSE - Extract command revision
                //-------------------------------------------------------------
                RX_PARSE_CMDREV: begin
                    $display("[CONTROLLER][RX_PARSE_CMDREV] cmd_pos 0x%02X, rx_byte 0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_CMDREV;
                    case (cmd_pos)
                        3'd0: begin
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            // Check REPORT byte
                            if (com_rx_byte == REPORT_NORMAL) begin
                                $display("[CONTROLLER][RX_PARSE_CMDREV] REPORT_NORMAL received");
                                com_rx_next <= 1'b1;     // Advance to revision data
                                main_state <= STATE_RX_NEXT;
                            end else begin
                                $display("[CONTROLLER][RX_PARSE_CMDREV] ERROR: Bad REPORT 0x%02X for CMDREV", com_rx_byte);
                                $display("[CONTROLLER][FATAL_ERROR] CMDREV failed - device cannot provide command revision");
                                main_state <= STATE_FATAL_ERROR;
                            end
                        end
                        3'd1: begin
                            // Store command revision (BCD format)
                            jvs_nodes_r.node_cmd_ver[current_device_addr - 1] <= com_rx_byte;
                            $display("[CONTROLLER][RX_PARSE_CMDREV] Command revision stored: 0x%02X", com_rx_byte);
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= CMDREV_TO_JVSREV_DELAY;
                            return_state <= STATE_SEND_JVSREV;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                            $display("[CONTROLLER] CMDREV complete, adding %0d cycle delay before JVSREV", CMDREV_TO_JVSREV_DELAY);
                        end
                        default: begin
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= CMDREV_TO_JVSREV_DELAY;
                            return_state <= STATE_SEND_JVSREV;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                        end
                    endcase
                end
                
                //-------------------------------------------------------------
                // JVS REVISION REQUEST - Get JVS protocol revision
                //-------------------------------------------------------------
                STATE_SEND_JVSREV: begin
                    // Send JVSREV command using sequential byte transmission
                    if (com_tx_ready) begin
                        com_dst_node <= current_device_addr; // 01
                        return_state <= STATE_SEND_JVSREV;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_JVSREV;          // Command revision command (0x11)
                                com_tx_cmd_push <= 1'b1;            // Push as command
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end
                end
                
                //-------------------------------------------------------------
                // PARSE JVSREV RESPONSE - Extract JVS revision
                //-------------------------------------------------------------
                RX_PARSE_JVSREV: begin
                    $display("[CONTROLLER][RX_PARSE_JVSREV] cmd_pos 0x%02X, rx_byte 0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_JVSREV;
                    case (cmd_pos)
                        3'd0: begin
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            // Check REPORT byte
                            if (com_rx_byte == REPORT_NORMAL) begin
                                $display("[CONTROLLER][RX_PARSE_JVSREV] REPORT_NORMAL received");
                                com_rx_next <= 1'b1;     // Advance to revision data
                                main_state <= STATE_RX_NEXT;
                            end else begin
                                $display("[CONTROLLER][RX_PARSE_JVSREV] ERROR: Bad REPORT 0x%02X for JVSREV", com_rx_byte);
                                $display("[CONTROLLER][FATAL_ERROR] JVSREV failed - device cannot provide JVS revision");
                                main_state <= STATE_FATAL_ERROR;
                            end
                        end
                        3'd1: begin
                            // Store JVS revision (BCD format)
                            jvs_nodes_r.node_jvs_ver[current_device_addr - 1] <= com_rx_byte;
                            $display("[CONTROLLER][RX_PARSE_JVSREV] JVS revision stored: 0x%02X", com_rx_byte);
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= JVSREV_TO_COMMVER_DELAY;
                            return_state <= STATE_SEND_COMMVER;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                            $display("[CONTROLLER] JVSREV complete, adding %0d cycle delay before COMMVER", JVSREV_TO_COMMVER_DELAY);
                        end
                        default: begin
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= JVSREV_TO_COMMVER_DELAY;
                            return_state <= STATE_SEND_COMMVER;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                        end
                    endcase
                end
                
                //-------------------------------------------------------------
                // COMMUNICATIONS VERSION REQUEST - Get communication version
                //-------------------------------------------------------------
                STATE_SEND_COMMVER: begin
                    // Send COMMVER command using sequential byte transmission
                    if (com_tx_ready) begin
                        // Initialize command parameters on first entry
                        com_dst_node <= current_device_addr; // 01
                        return_state <= STATE_SEND_COMMVER;
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_COMMVER;          // Command revision command (0x11)
                                com_tx_cmd_push <= 1'b1;            // Push as command
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end
                end
                
                //-------------------------------------------------------------
                // PARSE COMMVER RESPONSE - Extract communications version
                //-------------------------------------------------------------
                RX_PARSE_COMMVER: begin
                    $display("[CONTROLLER][RX_PARSE_COMMVER] cmd_pos 0x%02X, rx_byte 0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_COMMVER;
                    case (cmd_pos)
                        3'd0: begin
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            // Check REPORT byte
                            if (com_rx_byte == REPORT_NORMAL) begin
                                $display("[CONTROLLER][RX_PARSE_COMMVER] REPORT_NORMAL received");
                                com_rx_next <= 1'b1;     // Advance to revision data
                                main_state <= STATE_RX_NEXT;
                            end else begin
                                $display("[CONTROLLER][RX_PARSE_COMMVER] ERROR: Bad REPORT 0x%02X for COMMVER", com_rx_byte);
                                $display("[CONTROLLER][FATAL_ERROR] COMMVER failed - device cannot provide communications version");
                                main_state <= STATE_FATAL_ERROR;
                            end
                        end
                        3'd1: begin
                            // Store communications version (BCD format)
                            jvs_nodes_r.node_com_ver[current_device_addr - 1] <= com_rx_byte;
                            $display("[CONTROLLER][RX_PARSE_COMMVER] Communications version stored: 0x%02X", com_rx_byte);
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= COMMVER_TO_FEATURES_DELAY;
                            return_state <= STATE_SEND_FEATCHK;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                            $display("[CONTROLLER] COMMVER complete, adding %0d cycle delay before FEATCHK", COMMVER_TO_FEATURES_DELAY);
                        end
                        default: begin
                            cmd_pos <= 8'd0;          // Reset position for next command
                            delay_counter <= COMMVER_TO_FEATURES_DELAY;
                            return_state <= STATE_SEND_FEATCHK;
                            main_state <= STATE_MAIN_TIMER_DELAY;
                        end
                    endcase
                end
                
                //-------------------------------------------------------------
                // FEATURE CHECK REQUEST - Get device capabilities
                //-------------------------------------------------------------
                STATE_SEND_FEATCHK: begin
                    // Send FEATCHK command using sequential byte transmission
                    if (com_tx_ready) begin
                        // Initialize command parameters on first entry
                        if (cmd_pos == 0) begin
                            com_dst_node <= current_device_addr; // 01
                            return_state <= STATE_SEND_FEATCHK;
                        end
                        
                        // Select byte and signal based on position
                        case (cmd_pos)
                            3'd0: begin
                                com_tx_data <= CMD_FEATCHK;         // Feature check command (0x14)
                                com_tx_cmd_push <= 1'b1;            // Push as command
                                main_state <= STATE_TX_NEXT;        // Go to TX_NEXT
                            end
                            default: begin
                                // All bytes sent, commit and transition
                                com_commit <= 1'b1;
                                cmd_pos <= 8'd0;
                                main_state <= STATE_WAIT_RX;
                            end
                        endcase
                    end
                end

                RX_PARSE_FEATURES: begin
                    $display("[CONTROLLER][RX_PARSE_FEATURES] cmd_pos 0x%02X, rx_byte 0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_FEATURES;
                    case (cmd_pos)
                        3'd0: begin
                            // Check REPORT byte
                            com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                            if (com_rx_byte == REPORT_NORMAL) begin
                                $display("[CONTROLLER][FEATCHK] Report Normal");
                                com_rx_next <= 1'b1;
                                return_state <= RX_PARSE_FEATURES_FUNCS;
                                main_state <= STATE_RX_NEXT;
                                cmd_pos <= 0; // set cmd_pos to 0 for functions parsing, RX_NEXT increment cmd_pos so func parsing start a 1
                            end else begin
                                $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for COMMVER", com_rx_byte);
                                main_state <= STATE_WAIT_RX;
                            end
                        end
                    endcase
                end
                RX_PARSE_FEATURES_FUNCS: begin
                    $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] cmd_pos 0x%02X, rx_byte 0x%02X, rx_remaining=%d", cmd_pos, com_rx_byte, com_rx_remaining);
                    return_state <= RX_PARSE_FEATURES_FUNCS;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd1: begin // FUNC
                                if (com_rx_byte == 8'h00) begin
                                    // Terminator found - feature parsing complete
                                    $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Feature parsing complete (terminator found)");
                                    $display("[CONTROLLER] *** JVS INITIALIZATION COMPLETE - ACTIVATING jvs_data_ready_init ***");
                                    jvs_data_ready_init <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    // Add delay before going to input polling
                                    delay_counter <= FEATURES_TO_IDLE_DELAY;
                                    return_state <= STATE_SEND_INPUTS;
                                    main_state <= STATE_MAIN_TIMER_DELAY;
                                    $display("[CONTROLLER] FEATURES complete, adding %0d cycle delay before polling", FEATURES_TO_IDLE_DELAY);
                                end else begin
                                    // Store function code and continue
                                    current_func_code <= com_rx_byte;
                                    $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Parsing function 0x%02X", com_rx_byte);
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            3'd2: begin // ARG1
                                $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Parsing arg1 0x%02X for func 0x%02X", com_rx_byte, current_func_code);
                                case (current_func_code)
                                    FUNC_INPUT_DIGITAL: begin
                                        jvs_nodes_r.node_players[current_device_addr - 1] <= com_rx_byte[3:0];
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Digital: %d players", com_rx_byte[3:0]);
                                    end
                                    FUNC_INPUT_COIN: begin
                                        jvs_nodes_r.node_coin_slots[current_device_addr - 1] <= com_rx_byte[3:0];
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Coin: %d slots", com_rx_byte[3:0]);
                                    end
                                    FUNC_INPUT_ANALOG: begin
                                        jvs_nodes_r.node_analog_channels[current_device_addr - 1] <= com_rx_byte[3:0];
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Analog: %d channels", com_rx_byte[3:0]);
                                    end
                                    FUNC_INPUT_ROTARY: begin
                                        jvs_nodes_r.node_rotary_channels[current_device_addr - 1] <= com_rx_byte[3:0];
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Rotary: %d channels", com_rx_byte[3:0]);
                                    end
                                    FUNC_INPUT_KEYCODE: begin
                                        jvs_nodes_r.node_has_keycode_input[current_device_addr - 1] <= 1'b1;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Keycode input supported");
                                    end
                                    FUNC_INPUT_SCREEN_POS: begin
                                        jvs_nodes_r.node_screen_pos_x_bits[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Screen: %d X bits", com_rx_byte);
                                    end
                                    FUNC_INPUT_MISC_DIGITAL: begin
                                        jvs_nodes_r.node_misc_digital_inputs[current_device_addr - 1][15:8] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Misc digital: MSB=0x%02X", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_CARD: begin
                                        jvs_nodes_r.node_card_system_slots[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] %d Cards system present", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_HOPPER: begin
                                        jvs_nodes_r.node_medal_hopper_channels[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] %d Medal Hopper channels", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_DIGITAL: begin
                                        jvs_nodes_r.node_digital_outputs[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Digital outputs: %d channels", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_ANALOG: begin
                                        jvs_nodes_r.node_analog_output_channels[current_device_addr - 1] <= com_rx_byte[3:0];
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Analog outputs: %d channels", com_rx_byte[3:0]);
                                    end
                                    FUNC_OUTPUT_CHAR: begin
                                        jvs_nodes_r.node_has_char_display[current_device_addr - 1] <= 1'b1;
                                        jvs_nodes_r.node_char_display_width[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Character display: %d width", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_BACKUP: begin
                                        jvs_nodes_r.node_has_backup[current_device_addr - 1] <= 1'b1;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Backup present");
                                    end
                                    default: begin
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Unknown function 0x%02X, arg1=0x%02X", current_func_code, com_rx_byte);
                                    end
                                endcase
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            3'd3: begin // ARG2
                                $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Parsing arg2 0x%02X for func 0x%02X", com_rx_byte, current_func_code);
                                case (current_func_code)
                                    FUNC_INPUT_DIGITAL: begin
                                        jvs_nodes_r.node_buttons[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Digital: %d buttons per player", com_rx_byte);
                                    end
                                    FUNC_INPUT_ANALOG: begin
                                        jvs_nodes_r.node_analog_bits[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Analog: %d bits resolution", com_rx_byte);
                                    end
                                    FUNC_INPUT_SCREEN_POS: begin
                                        jvs_nodes_r.node_screen_pos_y_bits[current_device_addr - 1] <= com_rx_byte;
                                        jvs_nodes_r.node_has_screen_pos[current_device_addr - 1] <= 1'b1;
                                        has_screen_pos <= 1'b1;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Screen: %d Y bits", com_rx_byte);
                                    end
                                    FUNC_INPUT_MISC_DIGITAL: begin
                                        jvs_nodes_r.node_misc_digital_inputs[current_device_addr - 1][7:0] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Misc digital: LSB=0x%02X", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_CHAR: begin
                                        jvs_nodes_r.node_char_display_height[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Character display: %d height", com_rx_byte);
                                    end
                                    default: begin
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Function 0x%02X arg2=0x%02X (unused)", current_func_code, com_rx_byte);
                                    end
                                endcase
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            3'd4: begin // ARG3
                                $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Parsing arg3 0x%02X for func 0x%02X", com_rx_byte, current_func_code);
                                case (current_func_code)
                                    FUNC_INPUT_SCREEN_POS: begin
                                        jvs_nodes_r.node_screen_pos_channels[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Screen: %d channels", com_rx_byte);
                                    end
                                    FUNC_OUTPUT_CHAR: begin
                                        jvs_nodes_r.node_char_display_type[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Character display: type 0x%02X", com_rx_byte);
                                    end
                                    default: begin
                                        $display("[CONTROLLER][RX_PARSE_FEATURES_FUNCS] Function 0x%02X arg3=0x%02X (unused)", current_func_code, com_rx_byte);
                                    end
                                endcase
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                                cmd_pos <= 0; // end of FUNC ARGS
                            end
                        endcase
                    end else begin
                        main_state <= STATE_SEND_INPUTS;
                    end
                end

                //-------------------------------------------------------------
                // READ INPUTS COMMAND - Request current input states
                //-------------------------------------------------------------
                STATE_SEND_INPUTS: begin
                    // Send input commands using new jvs_com interface
                    if (com_tx_ready) begin
                        // Set destination node
                        com_dst_node <= current_device_addr; // 01

                        // Reset cmd_pos for new polling cycle
                        cmd_pos <= 8'd0;

                        // Begin progressive state machine - start with switch inputs
                        main_state <= STATE_SEND_INPUTS_SWITCH;
                    end
                end

                //-------------------------------------------------------------
                // INPUT BUILDING PROGRESSIVE STATES
                //-------------------------------------------------------------
                STATE_SEND_INPUTS_SWITCH: begin
                    if (jvs_nodes_r.node_players[current_device_addr - 1] > 0) begin
                        // Send SWINP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_SWITCH;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_SWINP;         // SWINP command (0x20)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= jvs_nodes_r.node_players[current_device_addr - 1];  // Number of players
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd2: begin
                                    com_tx_data <= (jvs_nodes_r.node_buttons[current_device_addr - 1] + 7) / 8; // Bytes for buttons
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_COIN;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_COIN;
                    end
                end
                STATE_SEND_INPUTS_COIN: begin // (CMD_COININP) @TODO: (CMD_COINDEC),(COININC)
                    if (jvs_nodes_r.node_coin_slots[current_device_addr - 1] > 0) begin
                        // Send COININP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_COIN;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_COININP;       // COININP command (0x21)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= jvs_nodes_r.node_coin_slots[current_device_addr - 1]; // Number of coin slots
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_ANALOG;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_ANALOG;
                    end
                end
                STATE_SEND_INPUTS_ANALOG: begin
                    if (jvs_nodes_r.node_analog_channels[current_device_addr - 1] > 0) begin
                        // Send ANLINP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_ANALOG;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_ANLINP;        // ANLINP command (0x22)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= jvs_nodes_r.node_analog_channels[current_device_addr - 1]; // Number of analog channels
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_ROTARY;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_ROTARY;
                    end
                end
                STATE_SEND_INPUTS_ROTARY: begin
                    if (jvs_nodes_r.node_rotary_channels[current_device_addr - 1] > 0) begin
                        // Send ROTINP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_ROTARY;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_ROTINP;        // ROTINP command (0x23)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= jvs_nodes_r.node_rotary_channels[current_device_addr - 1]; // Number of rotary channels
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_KEYCODE;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_KEYCODE;
                    end
                end
                STATE_SEND_INPUTS_KEYCODE: begin
                    if (jvs_nodes_r.node_has_keycode_input[current_device_addr - 1]) begin
                        // Send KEYINP command using sequential byte transmission (no parameters)
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_KEYCODE;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_KEYINP;        // KEYINP command (0x24)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_SCREEN;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_SCREEN;
                    end
                end
                STATE_SEND_INPUTS_SCREEN: begin
                    if (jvs_nodes_r.node_has_screen_pos[current_device_addr - 1]) begin
                        // Send SCRPOSINP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_SCREEN;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_SCRPOSINP;     // SCRPOSINP command (0x25)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= 8'h01;            // Channel index
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_INPUTS_MISC;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_INPUTS_MISC;
                    end
                end
                STATE_SEND_INPUTS_MISC: begin
                    if (jvs_nodes_r.node_misc_digital_inputs[current_device_addr - 1] > 0) begin
                        // Send MISCSWINP command using sequential byte transmission
                        if (com_tx_ready) begin
                            // Initialize command parameters on first entry
                            if (cmd_pos == 0) begin
                                com_dst_node <= current_device_addr;
                                return_state <= STATE_SEND_INPUTS_MISC;
                            end

                            // Select byte and signal based on position
                            case (cmd_pos)
                                3'd0: begin
                                    com_tx_data <= CMD_MISCSWINP;     // MISCSWINP command (0x26)
                                    com_tx_cmd_push <= 1'b1;         // Push as command
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                3'd1: begin
                                    com_tx_data <= (jvs_nodes_r.node_misc_digital_inputs[current_device_addr - 1] + 7) / 8; // Bytes needed
                                    com_tx_data_push <= 1'b1;        // Push as data
                                    main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                end
                                default: begin
                                    // All bytes sent, commit and transition
                                    //com_commit <= 1'b1;
                                    cmd_pos <= 8'd0;
                                    main_state <= STATE_SEND_OUTPUT_DIGITAL;
                                end
                            endcase
                        end
                    end else begin
                        main_state <= STATE_SEND_OUTPUT_DIGITAL;
                    end
                end
                // @TODO: Card system not supported
                // @TODO: Medal Hopper not supported (CMD_PAYCNT),(PAYINC),
                STATE_SEND_OUTPUT_DIGITAL: begin // (CMD_OUTPUT1) @TODO: (CMD_OUTPUT2),(CMD_OUTPUT3)
                    // Check if device has digital outputs
                    if (jvs_nodes_r.node_digital_outputs[current_device_addr - 1] > 0) begin
                        if (jvs_nodes_r.node_players[current_device_addr - 1] == 1) begin
                            // Single player mode (Time Crisis style) - Send OUTPUT1 command using sequential byte transmission
                            if (com_tx_ready) begin
                                // Initialize command parameters on first entry
                                if (cmd_pos == 0) begin
                                    com_dst_node <= current_device_addr;
                                    return_state <= STATE_SEND_OUTPUT_DIGITAL;
                                end

                                // Select byte and signal based on position
                                case (cmd_pos)
                                    3'd0: begin
                                        com_tx_data <= CMD_OUTPUT1;       // OUTPUT1 command (0x32)
                                        com_tx_cmd_push <= 1'b1;         // Push as command
                                        main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                    end
                                    3'd1: begin
                                        com_tx_data <= 8'h03;            // send 3 bytes
                                        com_tx_data_push <= 1'b1;        // Push as data
                                        main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                    end
                                    3'd2: begin
                                        com_tx_data <= gpio_output_value; // Set GPIO1 to current value from SNAC
                                        com_tx_data_push <= 1'b1;        // Push as data
                                        main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                    end
                                    3'd3: begin
                                        com_tx_data <= 8'hA0;            // do not know what A is for, but taken from TC4 capture
                                        com_tx_data_push <= 1'b1;        // Push as data
                                        main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                    end
                                    3'd4: begin
                                        com_tx_data <= 8'h00;
                                        com_tx_data_push <= 1'b1;        // Push as data
                                        main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                    end
                                    default: begin
                                        // All bytes sent, transition to finalize
                                        cmd_pos <= 8'd0;
                                        main_state <= STATE_SEND_OUTPUT_ANALOG;
                                        current_channel <= 8'd0;
                                    end
                                endcase
                            end
                        end else begin
                            cmd_pos <= 8'd0;
                            main_state <= STATE_SEND_OUTPUT_ANALOG;
                            current_channel <= 8'd0;
                        end
                    end else begin
                        cmd_pos <= 8'd0;
                        main_state <= STATE_SEND_OUTPUT_ANALOG;
                        current_channel <= 8'd0;
                    end
                end
                // @TODO: Analog Output not supported (CMD_ANLOUT)
                STATE_SEND_OUTPUT_ANALOG: begin // (CMD_ANLOUT)
                    // Check if device has analog outputs
                    if (jvs_nodes_r.node_analog_output_channels[current_device_addr - 1] > 0) begin
                        if(com_tx_ready) begin
                               // Initialize command parameters on first entry
                                if (cmd_pos == 0) begin
                                    com_dst_node <= current_device_addr;
                                    return_state <= STATE_SEND_OUTPUT_ANALOG;
                                end
                                if(current_channel >= jvs_nodes_r.node_analog_output_channels[current_device_addr - 1]) begin
                                    main_state <= STATE_SEND_FINALIZE;
                                    cmd_pos <= 0;
                                end else begin
                                    case (cmd_pos)
                                        3'd0: begin
                                            current_channel <= 0;
                                            com_tx_data <= CMD_ANLOUT;       // OUTPUT1 command (0x33)
                                            com_tx_cmd_push <= 1'b1;         // Push as command
                                            main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                        end
                                        3'd1: begin
                                            com_tx_data <= jvs_nodes_r.node_analog_output_channels[current_device_addr - 1]; // Number of channels to send
                                            com_tx_data_push <= 1'b1;
                                            main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                        end
                                        3'd2: begin
                                            com_tx_data <= 8'h00;           // Channel N MSB (@TODO: send null value at the momment)
                                            com_tx_data_push <=1'b1 ;       // Push data
                                            main_state <= STATE_TX_NEXT;    // Go to TX_NEXT
                                        end
                                        3'd3: begin
                                            com_tx_data <= 8'h00;            // Channel N LSB (@TODO: send null value at the momment)
                                            com_tx_data_push <= 1'b1;       // Push data
                                            main_state <= STATE_TX_NEXT;     // Go to TX_NEXT
                                            current_channel <= current_channel + 1;
                                            cmd_pos <= 1; // Go back to "3'd2" (MSB of next channel) after increased by TX_NEXT
                                        end
                                    endcase
                                end
                        end else begin
                            main_state <= STATE_SEND_FINALIZE;
                        end
                    end else begin
                        main_state <= STATE_SEND_FINALIZE;
                    end
                end
                /*
                Command name
                    Analog Outputs
                    byte0
                    byte1
                    byte2
                    byte3
                    ...
                    byteN
                    Request Data
                    33, channel, data, ...
                    33
                    Command Code
                    (02)
                    Channel count
                    (18)
                    Channel 1 MSB
                    (01)
                    Channel 1 LSB
                    ...
                    ...
                    (4A)
                    Last Channel LSB
                    Response Data
                    01 (report)
                    (01)
                    –
                    –
                    –
                    –
                    –
                    Report
                    Outputs data to analog outputs. Analog data is always specified as 16 bits, with the valid bits being
                    moved to the top, and the remainder set to 0. In this way, main board software does not need to know the
                    precision of the analog data.
                */
                // @TODO: Characters Output not supported (CHAROUT)
                // @TODO: Backup not support
                //-------------------------------------------------------------
                // FINALIZE MULTI-COMMAND FRAME - Commit all accumulated commands
                //-------------------------------------------------------------
                STATE_SEND_FINALIZE: begin
                    $display("[CONTROLLER][STATE_SEND_FINALIZE] Committing multi-command frame");
                    com_commit <= 1'b1;
                    cmd_pos <= 8'd0;
                    main_state <= STATE_WAIT_RX;
                end

                RX_PARSE_INPUT_CMD: begin
                    $display("[CONTROLLER][RX_PARSE_INPUT_CMD] Parsing command 0x%02X, cmd_pos=%d, rx_byte=0x%02X, cmd_count=%d", com_src_cmd, cmd_pos, com_rx_byte, com_src_cmd_count);
                    // Check if there are commands in the FIFO
                    if (com_src_cmd_count > 0 && com_rx_remaining > 0) begin
                        // Parse based on current command in FIFO
                        case (com_src_cmd)
                            CMD_SETADDR: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][SETADDR] Address %d accepted", current_device_addr);
                                            cmd_pos <= 8'd0;
                                            main_state <= STATE_SEND_IOIDENT;
                                        end else begin
                                            $display("[CONTROLLER][SETADDR] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                endcase
                            end
                            CMD_IOIDENT: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            copy_write_idx <= 8'd0;  // Reset write index for name copying
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][IOIDENT] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                    default: begin
                                        // Copy device name characters until null terminator or end of data
                                        if (com_rx_remaining > 0) begin
                                            if (com_rx_byte == 8'h00) begin
                                                // Found null terminator, store it and finish copying
                                                jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= 8'h00;
                                                $display("[CONTROLLER][IOIDENT] Name copy complete, %d chars", copy_write_idx);
                                                cmd_pos <= 8'd0;
                                                main_state <= STATE_SEND_CMDREV;
                                            end else if (copy_write_idx < jvs_node_info_pkg::NODE_NAME_SIZE - 1) begin
                                                // Store character and advance
                                                jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= com_rx_byte;
                                                copy_write_idx <= copy_write_idx + 1;
                                                return_state <= RX_PARSE_INPUT_CMD;
                                                main_state <= STATE_RX_NEXT;
                                                com_rx_next <= 1'b1;
                                            end else begin
                                                // Name too long, truncate and finish
                                                jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= 8'h00;
                                                $display("[CONTROLLER][IOIDENT] Name truncated at %d chars", copy_write_idx);
                                                cmd_pos <= 8'd0;
                                                main_state <= STATE_SEND_CMDREV;
                                            end
                                        end else begin
                                            // No more data, finish name copy
                                            jvs_nodes_r.node_name[current_device_addr - 1][copy_write_idx] <= 8'h00;
                                            cmd_pos <= 8'd0;
                                            main_state <= STATE_SEND_CMDREV;
                                        end
                                    end
                                endcase
                            end
                            CMD_CMDREV: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][CMDREV] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                    3'd1: begin
                                        // Store command revision (BCD format)
                                        jvs_nodes_r.node_cmd_ver[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][CMDREV] Command revision: 0x%02X", com_rx_byte);
                                        cmd_pos <= 8'd0;
                                        main_state <= STATE_SEND_JVSREV;
                                    end
                                endcase
                            end
                            CMD_JVSREV: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][JVSREV] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                    3'd1: begin
                                        // Store JVS revision (BCD format)
                                        jvs_nodes_r.node_jvs_ver[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][JVSREV] JVS revision: 0x%02X", com_rx_byte);
                                        cmd_pos <= 8'd0;
                                        main_state <= STATE_SEND_COMMVER;
                                    end
                                endcase
                            end
                            CMD_COMMVER: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][COMMVER] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                    3'd1: begin
                                        // Store communication version (BCD format)
                                        jvs_nodes_r.node_com_ver[current_device_addr - 1] <= com_rx_byte;
                                        $display("[CONTROLLER][COMMVER] Communication version: 0x%02X", com_rx_byte);
                                        cmd_pos <= 8'd0;
                                        main_state <= STATE_SEND_FEATCHK;
                                    end
                                endcase
                            end
                            CMD_FEATCHK: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        com_src_cmd_next <= 1'b1; // Flush FIFO to advance to next command
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][FEATCHK] ERROR: Bad REPORT 0x%02X", com_rx_byte);
                                            main_state <= STATE_FATAL_ERROR;
                                        end
                                    end
                                    default: begin
                                        // Dispatch to RX_PARSE_FEATURES for feature parsing
                                        cmd_pos <= 0;
                                        main_state <= RX_PARSE_FEATURES;
                                    end
                                endcase
                            end
                            default: begin
                                $display("[CONTROLLER] Unknown command 0x%02X, advancing to next", com_src_cmd);
                                com_src_cmd_next <= 1'b1;
                                cmd_pos <= 0;
                                return_state <= RX_PARSE_INPUT_CMD;
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            CMD_SWINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][RX_PARSE_INPUT_CMD][SWINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER][RX_PARSE_INPUT_CMD][SWINP] ERROR: Bad REPORT 0x%02X for SWINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            cmd_pos <= 0;
                                            com_rx_next <= 1'b1;
                                            //main_state <= STATE_RX_NEXT;
                                            main_state <= STATE_FATAL_ERROR; // for now we stop the simulation @TODO: proper error handeling
                                        end
                                    end
                                    3'd1: begin
                                        $display("[CONTROLLER][RX_PARSE_INPUT_CMD][SWINP] Consume System byte %02X for SWINP", com_rx_byte);
                                        current_player <= 4'd0; // initialise player idx
                                        return_state <= RX_PARSE_SWINP;
                                        cmd_pos <= 0;
                                        main_state <= STATE_RX_NEXT;
                                        com_rx_next <= 1'b1;
                                    end
                                endcase
                            end
                            CMD_COININP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][COININP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                            current_coin <= 0; // Initialize coin counter for parsing
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for COININP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            com_rx_next <= 1'b1;
                                            //main_state <= STATE_RX_NEXT;
                                            main_state <= STATE_FATAL_ERROR; // for now we stop the simulation @TODO: proper error handeling
                                        end
                                    end
                                    3'd1: begin
                                        // Dispatch to specialized ANLINP state
                                        $display("[CONTROLLER] Dispatching to ANLINP specialized parser");
                                        return_state <= RX_PARSE_COININP;
                                        main_state <= RX_PARSE_COININP;
                                    end
                                endcase
                            end
                            CMD_ANLINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][ANLINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for ANLINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    3'd1: begin
                                        // Dispatch to specialized ANLINP state
                                        $display("[CONTROLLER] Dispatching to ANLINP specialized parser");
                                        cmd_pos <= 0;
                                        return_state <= RX_PARSE_ANLINP;
                                        main_state <= RX_PARSE_ANLINP;
                                    end
                                endcase
                            end
                            CMD_ROTINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][ROTINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for ROTINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    default: begin
                                        // Simple parsing - skip rotary data (not implemented)
                                        $display("[CONTROLLER] Skipping ROTINP byte: 0x%02X", com_rx_byte);
                                        // Check if more data or advance to next command
                                        if (com_rx_remaining <= 1) begin
                                            // Last byte, advance to next command
                                            $display("[CONTROLLER] ROTINP parsing complete");
                                            cmd_pos <= 0;
                                            com_src_cmd_next <= 1'b1;
                                        end
                                        return_state <= RX_PARSE_INPUT_CMD;
                                        main_state <= STATE_RX_NEXT;
                                        com_rx_next <= 1'b1;
                                    end
                                endcase
                            end
                            CMD_KEYINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][KEYINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for KEYINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    default: begin
                                        // Simple parsing - skip keycode data (not implemented)
                                        $display("[CONTROLLER] Skipping KEYINP byte: 0x%02X", com_rx_byte);
                                        // Check if more data or advance to next command
                                        if (com_rx_remaining <= 1) begin
                                            // Last byte, advance to next command
                                            $display("[CONTROLLER] KEYINP parsing complete");
                                            cmd_pos <= 0;
                                            com_src_cmd_next <= 1'b1;
                                        end
                                        return_state <= RX_PARSE_INPUT_CMD;
                                        main_state <= STATE_RX_NEXT;
                                        com_rx_next <= 1'b1;
                                    end
                                endcase
                            end
                            CMD_SCRPOSINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][SCRPOSINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for SCRPOSINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    3'd1: begin
                                        // Dispatch to specialized SCRPOSINP state for screen position parsing
                                        $display("[CONTROLLER] Dispatching to SCRPOSINP specialized parser");
                                        cmd_pos <= 0;
                                        return_state <= RX_PARSE_SCRPOSINP;
                                        main_state <= RX_PARSE_SCRPOSINP;
                                    end
                                endcase
                            end
                            CMD_MISCSWINP: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][MISCSWINP] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for MISCSWINP", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    default: begin
                                        // Simple parsing - skip misc digital data (not implemented)
                                        $display("[CONTROLLER] Skipping MISCSWINP byte: 0x%02X", com_rx_byte);
                                        // Check if more data or advance to next command
                                        if (com_rx_remaining <= 1) begin
                                            // Last byte, advance to next command
                                            $display("[CONTROLLER] MISCSWINP parsing complete");
                                            cmd_pos <= 0;
                                            com_src_cmd_next <= 1'b1;
                                        end
                                        return_state <= RX_PARSE_INPUT_CMD;
                                        main_state <= STATE_RX_NEXT;
                                        com_rx_next <= 1'b1;
                                    end
                                endcase
                            end
                            CMD_OUTPUT1: begin
                                case(cmd_pos)
                                    3'd0: begin
                                        // Check REPORT byte
                                        if (com_rx_byte == REPORT_NORMAL) begin
                                            $display("[CONTROLLER][OUTPUT1] Report Normal");
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end else begin
                                            $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for OUTPUT1", com_rx_byte);
                                            com_src_cmd_next <= 1'b1;
                                            cmd_pos <= 0;
                                            return_state <= RX_PARSE_INPUT_CMD;
                                            main_state <= STATE_RX_NEXT;
                                            com_rx_next <= 1'b1;
                                        end
                                    end
                                    default: begin
                                        // Simple parsing - OUTPUT1 response is just acknowledgment, no complex data
                                        $display("[CONTROLLER] OUTPUT1 acknowledgment byte: 0x%02X", com_rx_byte);
                                        // Check if more data or advance to next command
                                        if (com_rx_remaining <= 1) begin
                                            // Last byte, advance to next command
                                            $display("[CONTROLLER] OUTPUT1 parsing complete");
                                            cmd_pos <= 0;
                                            com_src_cmd_next <= 1'b1;
                                        end
                                        return_state <= RX_PARSE_INPUT_CMD;
                                        main_state <= STATE_RX_NEXT;
                                        com_rx_next <= 1'b1;
                                    end
                                endcase
                            end
                        endcase
                    end else begin
                        // No more commands, input parsing complete
                        $display("[CONTROLLER] All input commands processed, adding delay before next polling cycle");
                        jvs_data_ready_joy <= 1'b1; // Signal that input data is ready for gaming
                        // Add delay between polling cycles to avoid overwhelming the bus
                        delay_counter <= POLLING_INTERVAL_DELAY;
                        return_state <= STATE_SEND_INPUTS;
                        main_state <= STATE_MAIN_TIMER_DELAY;
                        $display("[CONTROLLER] Polling cycle complete, adding %0d cycle delay before next cycle", POLLING_INTERVAL_DELAY);
                    end
                end
                
                RX_PARSE_SWINP: begin
                    $display("[CONTROLLER][RX_PARSE_SWINP] Player=%d, cmd_pos=%d, rx_byte=0x%02X", current_player, cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_SWINP;
                    case (current_player)
                        4'd0: begin // Player 1
                            if (cmd_pos == 1) begin
                                $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P1 byte 1");
                                // First player data byte
                                p1_btn_state[15] <= com_rx_byte[7];  // START
                                p1_btn_state[14] <= com_rx_byte[6];  // SELECT/SERVICE
                                p1_btn_state[0]  <= com_rx_byte[5];  // UP
                                p1_btn_state[1]  <= com_rx_byte[4];  // DOWN
                                p1_btn_state[2]  <= com_rx_byte[3];  // LEFT
                                p1_btn_state[3]  <= com_rx_byte[2];  // RIGHT
                                p1_btn_state[4]  <= com_rx_byte[1];  // A (push1)
                                p1_btn_state[5]  <= com_rx_byte[0];  // B (push2)

                                if (jvs_nodes_r.node_buttons[current_device_addr - 1] <= 8) begin
                                    // Only 1 byte per player, clear unused bits and advance to next player
                                    p1_btn_state[13:6] <= 8'b00000000;
                                    current_player <= current_player + 1;
                                    cmd_pos <= 0;
                                end
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end else if (cmd_pos == 2 && jvs_nodes_r.node_buttons[current_device_addr - 1] > 8) begin
                                $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P1 byte 2");
                                // Second player data byte (additional buttons)
                                p1_btn_state[6] <= com_rx_byte[7];   // X (push3)
                                p1_btn_state[7] <= com_rx_byte[6];   // Y (push4)
                                p1_btn_state[8] <= com_rx_byte[5];   // push5 -> L1
                                p1_btn_state[9] <= com_rx_byte[4];   // push6 -> R1
                                p1_btn_state[10] <= com_rx_byte[3];  // push7 -> L2
                                p1_btn_state[11] <= com_rx_byte[2];  // push8 -> R2
                                p1_btn_state[12] <= com_rx_byte[1];  // push9 -> L3
                                p1_btn_state[13] <= com_rx_byte[0];  // push10 -> R3
                                // Advance to next player
                                current_player <= current_player + 1;
                                cmd_pos <= 0; // Reset for next player
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        end

                        4'd1: begin // Player 2
                            if (cmd_pos == 1) begin
                                $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P2 byte 1");
                                // First player data byte
                                p2_btn_state[15] <= com_rx_byte[7];  // START
                                p2_btn_state[14] <= com_rx_byte[6];  // SELECT/SERVICE
                                p2_btn_state[0]  <= com_rx_byte[5];  // UP
                                p2_btn_state[1]  <= com_rx_byte[4];  // DOWN
                                p2_btn_state[2]  <= com_rx_byte[3];  // LEFT
                                p2_btn_state[3]  <= com_rx_byte[2];  // RIGHT
                                p2_btn_state[4]  <= com_rx_byte[1];  // A (push1)
                                p2_btn_state[5]  <= com_rx_byte[0];  // B (push2)

                                if (jvs_nodes_r.node_buttons[current_device_addr - 1] <= 8) begin
                                    // Only 1 byte per player, clear unused bits and advance to next player
                                    p2_btn_state[13:6] <= 8'b00000000;
                                    current_player <= current_player + 1;
                                    cmd_pos <= 0;
                                end
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end else if (cmd_pos == 2 && jvs_nodes_r.node_buttons[current_device_addr - 1] > 8) begin
                                $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P2 byte 2");
                                // Second player data byte (additional buttons) - match your reference bit mapping
                                p2_btn_state[6] <= com_rx_byte[7];   // X (push3)
                                p2_btn_state[7] <= com_rx_byte[6];   // Y (push4)
                                p2_btn_state[8] <= com_rx_byte[5];   // push5 -> L1
                                p2_btn_state[9] <= com_rx_byte[4];   // push6 -> R1
                                p2_btn_state[10] <= com_rx_byte[3];  // push7 -> L2
                                p2_btn_state[11] <= com_rx_byte[2];  // push8 -> R2
                                // Clear unused upper bits for consistency with reference
                                p2_btn_state[13:12] <= 2'b00;
                                // Advance to next player
                                current_player <= current_player + 1;
                                cmd_pos <= 0; // Reset for next player
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        end

                        default: begin
                            if (current_player >= jvs_nodes_r.node_players[current_device_addr - 1]) begin
                                $display("[CONTROLLER][RX_PARSE_SWINP] All players processed, advancing to next command");
                                cmd_pos <= 0;
                                com_src_cmd_next <= 1'b1;
                                return_state <= RX_PARSE_INPUT_CMD;
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end else begin
                                // Additional players (if supported)
                                $display("[CONTROLLER][RX_PARSE_SWINP] Skipping unsupported player %d", current_player);
                                if (cmd_pos == 1) begin
                                    $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P%d byte 1", current_player);
                                    if (jvs_nodes_r.node_buttons[current_device_addr - 1] <= 8) begin
                                        // Only 1 byte per player, clear unused bits and advance to next player
                                        current_player <= current_player + 1;
                                        cmd_pos <= 0;
                                    end
                                    main_state <= STATE_FATAL_ERROR;
                                    com_rx_next <= 1'b1;
                                end
                                if (cmd_pos == 2 && jvs_nodes_r.node_buttons[current_device_addr - 1] > 8) begin
                                    $display("[CONTROLLER][RX_PARSE_SWINP] Parsing P%d byte 2", current_player);
                                    // Advance to next player
                                    current_player <= current_player + 1;
                                    cmd_pos <= 0; // Reset for next player
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                        end
                    endcase
                end

                RX_PARSE_COININP: begin
                    $display("[CONTROLLER][RX_PARSE_COININP] Parsing coin data, cmd_pos=%d, rx_byte=0x%02X, current_coin=%d", cmd_pos, com_rx_byte, current_coin);
                    if (com_rx_remaining > 0) begin
                        // Parse coin data (2 bytes per coin slot)
                        case (cmd_pos)
                            3'd1: begin // Parse byte 1 of current coin slot
                                // Format: [condition(2 bits) counter_MSB(6 bits)]
                                temp_coin_condition <= com_rx_byte[7:6];  // Top 2 bits = condition
                                temp_counter_msb <= com_rx_byte[5:0];     // Bottom 6 bits = counter MSB
                                $display("[CONTROLLER] Coin slot %d: condition=%d, msb=0x%02X", current_coin, com_rx_byte[7:6], com_rx_byte[5:0]);
                                return_state <= RX_PARSE_COININP;
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            3'd2: begin // Parse byte 2 of current coin slot then jump to next slot if needed
                                // Store complete coin data for this slot
                                coin_count[current_coin] <= {temp_counter_msb, com_rx_byte}; // 14-bit counter stored in 16-bit
                                
                                // Set coin increase signals based on condition (10 = increase)
                                case (current_coin)
                                    0: coin1 <= (temp_coin_condition == 2'b10);
                                    1: coin2 <= (temp_coin_condition == 2'b10);
                                    2: coin3 <= (temp_coin_condition == 2'b10);
                                    3: coin4 <= (temp_coin_condition == 2'b10);
                                endcase
                                
                                $display("[CONTROLLER] Coin slot %d: lsb=0x%02X, total=%d, increase=%b", 
                                        current_coin, com_rx_byte, {temp_counter_msb, com_rx_byte}, (temp_coin_condition == 2'b10));
                                
                                // Check if we need to parse the next coin slot
                                if (current_coin >= (jvs_nodes_r.node_coin_slots[current_device_addr - 1] - 1)) begin
                                    // Coin parsing complete, advance to next command
                                    $display("[CONTROLLER] Coin parsing complete, advancing to next command");
                                    cmd_pos <= 0;
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end else begin
                                    // Parse next coin slot
                                    current_coin <= current_coin + 1;
                                    cmd_pos <= 0; // Reset to parse next coin's first byte
                                    return_state <= RX_PARSE_COININP;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                        endcase
                    end else begin
                        // No more data, return to command dispatcher
                        cmd_pos <= 0;
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= return_state;
                    end
                end

                RX_PARSE_ANLINP: begin
                    $display("[CONTROLLER][RX_PARSE_ANLINP] Parsing analog data, cmd_pos=%d, rx_byte=0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_ANLINP;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd0: begin
                                // Check REPORT byte
                                if (com_rx_byte == REPORT_NORMAL) begin
                                    $display("[CONTROLLER][RX_PARSE_ANLINP] Report Normal");
                                    com_rx_next <= 1'b1;
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for ANLINP", com_rx_byte);
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            default: begin
                                // Parse analog input data based on node configuration
                                automatic logic [7:0] data_pos = cmd_pos - 1; // Adjust for REPORT byte
                                if (data_pos < (jvs_nodes_r.node_analog_channels[current_device_addr - 1] * 2)) begin // 2 bytes per channel
                                    automatic logic [3:0] channel_idx = data_pos / 2;
                                    if (data_pos % 2 == 0) begin
                                // High byte
                                case (channel_idx)
                                    0: p1_joy_state[31:24] <= com_rx_byte;  // P1 X axis high
                                    1: p1_joy_state[15:8] <= com_rx_byte;   // P1 Y axis high
                                    2: p2_joy_state[31:24] <= com_rx_byte;  // P2 X axis high
                                    3: p2_joy_state[15:8] <= com_rx_byte;   // P2 Y axis high
                                    default: begin
                                        // Store in screen position for channels > 3
                                        if (channel_idx == 4) screen_pos_x[15:8] <= com_rx_byte;
                                        else if (channel_idx == 5) screen_pos_y[15:8] <= com_rx_byte;
                                    end
                                endcase
                                $display("[CONTROLLER] Analog channel %d high byte: 0x%02X", channel_idx, com_rx_byte);
                            end else begin
                                // Low byte
                                case (channel_idx)
                                    0: p1_joy_state[23:16] <= com_rx_byte;  // P1 X axis low
                                    1: p1_joy_state[7:0] <= com_rx_byte;    // P1 Y axis low
                                    2: p2_joy_state[23:16] <= com_rx_byte;  // P2 X axis low
                                    3: p2_joy_state[7:0] <= com_rx_byte;    // P2 Y axis low
                                    default: begin
                                        // Store in screen position for channels > 3
                                        if (channel_idx == 4) screen_pos_x[7:0] <= com_rx_byte;
                                        else if (channel_idx == 5) screen_pos_y[7:0] <= com_rx_byte;
                                    end
                                endcase
                                $display("[CONTROLLER] Analog channel %d low byte: 0x%02X", channel_idx, com_rx_byte);
                            end
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end else begin
                                    // Analog parsing complete, check if more commands or return to polling
                                    $display("[CONTROLLER] Analog parsing complete, checking for more commands");
                                    cmd_pos <= 0;
                                    com_src_cmd_next <= 1'b1; // Advance to next command in FIFO
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                        endcase
                    end else begin
                        main_state <= STATE_IDLE;
                    end
                end

                //-------------------------------------------------------------
                // ADDITIONAL INPUT PARSING STATES - Not yet implemented
                //-------------------------------------------------------------
                RX_PARSE_ROTINP: begin
                    $display("[CONTROLLER][RX_PARSE_ROTINP] Parsing rotary data - pas encore implémenté");
                    return_state <= RX_PARSE_ROTINP;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd0: begin
                                // Check REPORT byte
                                if (com_rx_byte == REPORT_NORMAL) begin
                                    $display("[CONTROLLER][RX_PARSE_ROTINP] Report Normal");
                                    com_rx_next <= 1'b1;
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for ROTINP", com_rx_byte);
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            default: begin
                                // Parse rotary data - not yet implemented
                                $display("[CONTROLLER] Skipping rotary byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        endcase
                    end else begin
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= STATE_RX_NEXT;
                        com_rx_next <= 1'b1;
                    end
                end

                RX_PARSE_KEYINP: begin
                    $display("[CONTROLLER][RX_PARSE_KEYINP] Parsing keycode data - pas encore implémenté");
                    return_state <= RX_PARSE_KEYINP;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd0: begin
                                // Check REPORT byte
                                if (com_rx_byte == REPORT_NORMAL) begin
                                    $display("[CONTROLLER][RX_PARSE_KEYINP] Report Normal");
                                    com_rx_next <= 1'b1;
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for KEYINP", com_rx_byte);
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            default: begin
                                // Parse keycode data - not yet implemented
                                $display("[CONTROLLER] Skipping keycode byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        endcase
                    end else begin
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= STATE_RX_NEXT;
                        com_rx_next <= 1'b1;
                    end
                end

                RX_PARSE_SCRPOSINP: begin
                    $display("[CONTROLLER][RX_PARSE_SCRPOSINP] Parsing screen position data, cmd_pos=%d, rx_byte=0x%02X", cmd_pos, com_rx_byte);
                    return_state <= RX_PARSE_SCRPOSINP;
                    if (com_rx_remaining > 0) begin
                        // Parse screen position data (4 bytes: X_HIGH, X_LOW, Y_HIGH, Y_LOW)
                        // REPORT byte already consumed by RX_PARSE_INPUT_CMD, start parsing from cmd_pos=1
                        automatic logic [7:0] data_pos = cmd_pos - 1; // Adjust for REPORT byte
                        case (data_pos)
                            8'd0: begin // X coordinate high byte
                                screen_pos_x[15:8] <= com_rx_byte;
                                $display("[CONTROLLER] Screen X high byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            8'd1: begin // X coordinate low byte
                                screen_pos_x[7:0] <= com_rx_byte;
                                $display("[CONTROLLER] Screen X low byte: 0x%02X, X = %d", com_rx_byte, {screen_pos_x[15:8], com_rx_byte});
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            8'd2: begin // Y coordinate high byte
                                screen_pos_y[15:8] <= com_rx_byte;
                                $display("[CONTROLLER] Screen Y high byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            8'd3: begin // Y coordinate low byte
                                screen_pos_y[7:0] <= com_rx_byte;
                                $display("[CONTROLLER] Screen Y low byte: 0x%02X, Y = %d", com_rx_byte, {screen_pos_y[15:8], com_rx_byte});
                                $display("[CONTROLLER] Screen position complete: (%d, %d)", {screen_pos_x[15:8], screen_pos_x[7:0]}, {screen_pos_y[15:8], com_rx_byte});
                                // Screen position parsing complete, advance to next command
                                cmd_pos <= 0;
                                com_src_cmd_next <= 1'b1;
                                return_state <= RX_PARSE_INPUT_CMD;
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                            default: begin
                                // Unexpected data, skip
                                $display("[CONTROLLER] Unexpected SCRPOSINP data at pos %d: 0x%02X", data_pos, com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        endcase
                    end else begin
                        // No more data, return to command dispatcher
                        cmd_pos <= 0;
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= STATE_RX_NEXT;
                        com_rx_next <= 1'b1;
                    end
                end

                RX_PARSE_MISCSWINP: begin
                    $display("[CONTROLLER][RX_PARSE_MISCSWINP] Parsing misc digital data - pas encore implémenté");
                    return_state <= RX_PARSE_MISCSWINP;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd0: begin
                                // Check REPORT byte
                                if (com_rx_byte == REPORT_NORMAL) begin
                                    $display("[CONTROLLER][RX_PARSE_MISCSWINP] Report Normal");
                                    com_rx_next <= 1'b1;
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for MISCSWINP", com_rx_byte);
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            default: begin
                                // Parse misc digital data - not yet implemented
                                $display("[CONTROLLER] Skipping misc digital byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        endcase
                    end else begin
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= STATE_RX_NEXT;
                        com_rx_next <= 1'b1;
                    end
                end

                RX_PARSE_OUTPUT1: begin
                    $display("[CONTROLLER][RX_PARSE_OUTPUT1] Parsing output digital response - pas encore implémenté");
                    return_state <= RX_PARSE_OUTPUT1;
                    if (com_rx_remaining > 0) begin
                        case (cmd_pos)
                            3'd0: begin
                                // Check REPORT byte
                                if (com_rx_byte == REPORT_NORMAL) begin
                                    $display("[CONTROLLER][RX_PARSE_OUTPUT1] Report Normal");
                                    com_rx_next <= 1'b1;
                                    main_state <= STATE_RX_NEXT;
                                end else begin
                                    $display("[CONTROLLER] ERROR: Bad REPORT 0x%02X for OUTPUT1", com_rx_byte);
                                    com_src_cmd_next <= 1'b1;
                                    return_state <= RX_PARSE_INPUT_CMD;
                                    main_state <= STATE_RX_NEXT;
                                    com_rx_next <= 1'b1;
                                end
                            end
                            default: begin
                                // Parse output digital response - not yet implemented
                                $display("[CONTROLLER] Skipping output digital byte: 0x%02X", com_rx_byte);
                                main_state <= STATE_RX_NEXT;
                                com_rx_next <= 1'b1;
                            end
                        endcase
                    end else begin
                        com_src_cmd_next <= 1'b1;
                        return_state <= RX_PARSE_INPUT_CMD;
                        main_state <= STATE_RX_NEXT;
                        com_rx_next <= 1'b1;
                    end
                end

                //-------------------------------------------------------------
                // WAIT FOR DEVICE RESPONSE - Using edge detection for proper timing
                //-------------------------------------------------------------
                STATE_WAIT_RX: begin
                    if (com_rx_complete_negedge) begin
                        // Check STATUS byte decoded by jvs_com from received frame
                        if (com_src_cmd_status == STATUS_NORMAL) begin
                            // STATUS OK, dispatch to appropriate parser
                            $display("[CONTROLLER] PROCESSING 0x%02X with STATUS %02X", com_src_cmd, com_rx_byte);
                            cmd_pos <= 8'd0;
                            case (com_src_cmd)
                                CMD_SETADDR: main_state <= RX_PARSE_SETADDR;
                                CMD_IOIDENT: main_state <= RX_PARSE_IOIDENT;
                                CMD_CMDREV: main_state <= RX_PARSE_CMDREV;
                                CMD_JVSREV: main_state <= RX_PARSE_JVSREV;
                                CMD_COMMVER: main_state <= RX_PARSE_COMMVER;
                                CMD_FEATCHK: main_state <= RX_PARSE_FEATURES;
                                default: main_state <= RX_PARSE_INPUT_CMD; // For other commands, use unified parser
                            endcase
                        end else begin
                            // STATUS error, log and retry
                            $display("[CONTROLLER] ERROR: Bad STATUS 0x%02X for cmd 0x%02X", com_src_cmd_status, com_src_cmd);
                            case (com_src_cmd)
                                CMD_SETADDR: main_state <= STATE_FIRST_RESET;    // Critical - restart sequence
                                CMD_IOIDENT: main_state <= STATE_SEND_IOIDENT;     // Retry ID read
                                CMD_CMDREV: main_state <= STATE_SEND_CMDREV;     // Retry command revision
                                CMD_JVSREV: main_state <= STATE_SEND_JVSREV;     // Retry JVS revision
                                CMD_COMMVER: main_state <= STATE_SEND_COMMVER;   // Retry comm version
                                CMD_FEATCHK: main_state <= STATE_SEND_FEATCHK;   // Retry feature check
                                default: main_state <= STATE_IDLE;               // Continue with polling
                            endcase
                        end
                    //end else if (timeout_counter < 32'h0C3500) begin  // 10ms timeout - fast for responsive gaming
                    end else if (timeout_counter < RX_TIMEOUT_COUNT) begin  // 10ms timeout - fast for responsive gaming
                        timeout_counter <= timeout_counter + 1;
                    end else begin
                        $display("[CONTROLLER] RX_IDLE Timeout");
                        // Timeout handling - different strategies for different commands
                        case (com_src_cmd)
                            /*
                            CMD_SETADDR: main_state <= STATE_FIRST_RESET;    // Critical - restart sequence
                            CMD_IOIDENT: main_state <= STATE_SEND_IOIDENT;     // Retry ID read
                            CMD_CMDREV: main_state <= STATE_SEND_CMDREV;     // Retry command revision
                            CMD_JVSREV: main_state <= STATE_SEND_JVSREV;     // Retry JVS revision
                            CMD_COMMVER: main_state <= STATE_SEND_COMMVER;   // Retry comm version
                            CMD_FEATCHK: main_state <= STATE_SEND_FEATCHK;   // Retry feature check
                            */
                            default: main_state <= STATE_FATAL_ERROR;               // Continue with polling
                        endcase
                    end
                end

                //-------------------------------------------------------------
                // GENERIC TIMER DELAY STATE - Reusable delay for any state transition
                //-------------------------------------------------------------
                STATE_MAIN_TIMER_DELAY: begin
                    if (delay_counter > 0) begin
                        delay_counter <= delay_counter - 1;
                    end else begin
                        // Timer expired, return to caller state
                        main_state <= return_state;
                        $display("[CONTROLLER] MAIN_TIMER_DELAY complete, returning to state 0x%02X", return_state);
                    end
                end

                //-------------------------------------------------------------
                // GENERIC TX NEXT STATE - Handles pulse cleanup and position increment
                //-------------------------------------------------------------
                STATE_TX_NEXT: begin
                    $display("[CONTROLLER][STATE_TX_NEXT] cmd:%b data:%b commit:%b", com_tx_cmd_push, com_tx_data_push, com_commit);
                    $display("[CONTROLLER] STATE_TX_NEXT: clearing com_tx_cmd_push and com_tx_data_push");
                    com_tx_cmd_push <= 1'b0;
                    com_tx_data_push <= 1'b0;
                    cmd_pos <= cmd_pos + 1;
                    if(com_commit == 1'b1) begin
                        // Keep com_commit high until JVS_COM accepts it (tx_ready goes low)
                        if(!com_tx_ready) begin
                            // JVS_COM has accepted the commit (tx_ready went low)
                            com_commit <= 1'b0;
                            cmd_pos <= 8'h00;
                            main_state <= STATE_WAIT_RX;
                        end
                        // else: keep com_commit high and stay in TX_NEXT until JVS_COM is ready
                    end else begin
                        main_state <= return_state;
                    end
                end
                STATE_RX_NEXT: begin
                    $display("[CONTROLLER][STATE_RX_NEXT]");
                    com_rx_next <= 0;
                    cmd_pos <= cmd_pos + 1;                    
                    main_state <= return_state;
                end

                //-------------------------------------------------------------
                // FATAL ERROR STATE - Stop execution and display error
                //-------------------------------------------------------------
                STATE_FATAL_ERROR: begin
                    // Stay in error state and continuously display error message
                    $display("[CONTROLLER][FATAL_ERROR] JVS Controller has entered fatal error state");
                    $display("[CONTROLLER][FATAL_ERROR] System stopped for debugging");
                    
                    // Display jvs_nodes_r content for debugging
                    $display("[CONTROLLER][FATAL_ERROR] === JVS_NODES_R STATE DUMP ===");
                    for (int dev = 0; dev < 2; dev++) begin
                        $display("[FATAL_ERROR] Device %d:", dev);
                        $display("  node_id: 0x%02X", jvs_nodes_r.node_id[dev]);
                        $display("  node_cmd_ver: 0x%02X", jvs_nodes_r.node_cmd_ver[dev]);
                        $display("  node_jvs_ver: 0x%02X", jvs_nodes_r.node_jvs_ver[dev]);
                        $display("  node_com_ver: 0x%02X", jvs_nodes_r.node_com_ver[dev]);
                        $display("  node_players: %d", jvs_nodes_r.node_players[dev]);
                        $display("  node_buttons: %d", jvs_nodes_r.node_buttons[dev]);
                        $display("  node_analog_channels: %d", jvs_nodes_r.node_analog_channels[dev]);
                        $display("  node_analog_bits: %d", jvs_nodes_r.node_analog_bits[dev]);
                        $display("  node_coin_slots: %d", jvs_nodes_r.node_coin_slots[dev]);
                        $display("  node_rotary_channels: %d", jvs_nodes_r.node_rotary_channels[dev]);
                        $display("  node_digital_outputs: %d", jvs_nodes_r.node_digital_outputs[dev]);
                        $display("  node_analog_output_channels: %d", jvs_nodes_r.node_analog_output_channels[dev]);
                        $display("  node_has_keycode_input: %b", jvs_nodes_r.node_has_keycode_input[dev]);
                        $display("  node_has_screen_pos: %b", jvs_nodes_r.node_has_screen_pos[dev]);
                        if (jvs_nodes_r.node_has_screen_pos[dev]) begin
                            $display("    screen_pos_x_bits: %d", jvs_nodes_r.node_screen_pos_x_bits[dev]);
                            $display("    screen_pos_y_bits: %d", jvs_nodes_r.node_screen_pos_y_bits[dev]);
                        end
                        $display("  node_misc_digital_inputs: 0x%04X", jvs_nodes_r.node_misc_digital_inputs[dev]);
                        $display("  node_has_char_display: %b", jvs_nodes_r.node_has_char_display[dev]);
                        if (jvs_nodes_r.node_has_char_display[dev]) begin
                            $display("    char_display_width: %d", jvs_nodes_r.node_char_display_width[dev]);
                            $display("    char_display_height: %d", jvs_nodes_r.node_char_display_height[dev]);
                            $display("    char_display_type: 0x%02X", jvs_nodes_r.node_char_display_type[dev]);
                        end
                        $display("  node_has_backup: %b", jvs_nodes_r.node_has_backup[dev]);
                        
                        // Display device name
                        $write("  device_name: \"");
                        for (int i = 0; i < jvs_node_info_pkg::NODE_NAME_SIZE; i++) begin
                            if (jvs_nodes_r.node_name[dev][i] == 8'h00) break;
                            $write("%c", jvs_nodes_r.node_name[dev][i]);
                        end
                        $display("\"");
                    end
                    $display("[CONTROLLER][FATAL_ERROR] === END JVS_NODES_R DUMP ===");
                    
                    $finish; // Stop simulation immediately for debugging
                end

                //-------------------------------------------------------------
                // DEFAULT - Unknown state, go to fatal error
                //-------------------------------------------------------------
                default: begin
                    $display("[CONTROLLER][FATAL_ERROR] Unknown state 0x%02X - entering fatal error state", main_state);
                    main_state <= STATE_FATAL_ERROR;
                end
            endcase
        end
    end

endmodule